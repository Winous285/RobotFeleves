��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�   � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d PPINFwOEQ/ ��L A �!�%/� H� �&�)EQUIP 2� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CESS0s!_81s!J3�> �! � �$SOFT�T_�IDk2TOTAL7_EQs $�0�0�NO�2U SPI_OINDE]�5Xk2SCREEN_(4�_2SIGE0�_?q;�0PK_FI�� 	$THK�YGPANE�4 �� DUMMY1"dDDd!OE4LA!�R�!R�	 � �$TIT�!$I��N �Dd�Dd ��Dc@�D5�F6�F7*�F8�F9�G0�G�G@JA�E�GbA�E�G1�G� �F�G1�G2�B\�S�ASBN_C�F>"
 8F CN�V_J� ; �"�!_�CMNT�$F�LAGS]�CH�EC�8 � ELL�SETUP ރ $HO30IO��0� %�SMAC{RO�RREPR�X� D+�0��R{�T� UTOBACK�U�0 ��)DEVIC�CT	I*0�� �0�#��`B�S$INTE�RVALO#ISP�_UNI�O`_D�O>f7uiFR_F�0AIN�1���1<c�C_WAkda^�jOFF_O0N�DEL�hL� ?aA�a1b?9a�`C#?��P�1E��#s�ATB�d��MO<� �cE D [�M�c��^qREV��BILrw!XI�� QrR  �� OD�P�q$NO^PM�Wp�t�r/"�w� �u��q �p�0D`S� p E RD�_E�pCq$FS�SBn&$CHKBoD_SE^eAG �G�"$SLOT!_��2=�� V�d�%���3 a_ED�Im   � )�"��PS�`(4�%$EP�1�1$�OP�0�2�a�p_�OK�UST1P_�C� ��d��U �PLACI4!�Q�4�<( raCOMM� ,0$D����0�`���EOWBn�IGALL;OW� (K�":(2�0VARa��@h�2ao�L�0OUy�� ,Kvay��PS�`�0M_O]�����CF�t XF� GRP0��M=q�NFLI�ܓ�0U�IRE��$g"� S�WITCHړAX�_N�PSs"CF_��G� �� WARNM�`#!�!��qPLI�I�NST�� COR-0bF�LTRC�TRAT�PTE�� $AC�C1a�N ��r$�ORI�o"��RT��P_SFg CHUG�0I��rTא�1�I��T�I1�|�� x i#��Q��HDRBJ�; C,�2'�3'�4�'�5'�6'�7'�8�'�9s!ӡO`T <F П����#92^��LLECy�"MULTI�b�"N���1�!���0T_}R � 4F STY �"�R`�=l�)2`�p����`T |� @�&$c�Z`�pb��Pf�MO�0�TTOӰ:�Ew�EXT����pÁB���"2� ,��[0]�}Rദ�b�}�  D"}����Q���Q�kc	G���^ȇ1���ÂM���P�� 8ŋ� L�  ����P��`A��$J�OBn�/�i�G�TR;IG�  d�p�� ����³�7������!CO_M�b!� t�pF� CNG AiBA� ����M� ��!���p� �q��0���P[`��i�*�"6���0tB񉠎"MJ��_Rz�gC�QJ��$�?�Jk�D�%�C_�;������0ФR>�t#� �������G���0NHA;NC̳$LGa���B^a��� �D��A�`��gzRɡ�!�0�p�DB�3RA�AZ�0K�ELT�Ė��PFCT&��F�0�P��SM��cI��1� % ��% ��R��a����� S��&���M` 00{o e#HK~օA^S�������If_T$�"6SW�OCSXC)�?!%�h�p)3��T�$@�ΙPANN&�AIMG_HEIGHCr·WIDI AVT��0��H F_ASqPװ��`EXP�1|���CUST��U��&��|E\�%�C1NV _�`�a���' \%1y�`OR@�c,"�0gsk��PO��LBSYI�G��aR%��`좔Pspm��0k�DBPXWORK���(��$SKP_d�`ma�"<qTRp ) ���P��0�� �0�DJ!d/��_CN��R�#� �'PAL�S�Q�d�s�DKA7WAw'�^A�@�NFZpfBDBU��*L�"!PRS�7�
�8�Q����+ [pr�$1�$Z,
K�Li9,v?Ϣ�ʠR��-�?�4C��.�?ή4ENEy��� 1/�?�3J0RE`��2�0H��CuR+$L,C,$i3
�? �=KINE@�K!_D�I�RO�`�����ȳqvC��h �FPA4Ã3uR�PRN�B��MR��U!�u�CR�[@EWM �SIGN��A� .q�E��Q-$P��.3$Pp 2�/ P7�!PT2�PDu`L����VDBAR@�GO_AW���Jp �� �DCS�pZ�CYO_ 1���@1<�\�Q?fIG2�Z2>fN>�����
�qS&c}P�2 P $��R)B?�e�P=hPwg�Q#BYl�`gT+1�T/HNDG�23��KS��SE|�Q��SBL@㸣cc�T�qSL�4 HpZ ���V�TOFB�l�FE@fA�ǿb�TqSW5�b�DOC���MCS@�f�`Z$r�b H� �W0��T��rRSLA�V�16�rINP���f��LyqQP�7� $,�S���=�`�v��uFI��r줭sc�!��!9W1ԭrNTV'��r�V	��uSKIvT�E�@W���:�J�_� _�00�SAsFE�A�_SV��EXCLU��B J�PDJ L1�k�Y�d8�ƻrI_V� !�PPLY 0b���D9E~w��_ML2�B $VRFY_�#��Mk�IOU��憐� 0���:�O�P��L1S�@jb;�3572��Sr�� Px%X�{Pp�hs� �� 8 @Ɠ TA� qঠ {�c_SGN��96����@�A������iPt!��s"��~UN�0jdՔ�U���B �@� ��� �����!l�OGI�2:� @�`Fؒ���O�T�@@�:41(�774�C2�M`NI�2;��R������A�q��D{AY1#LOAD�T�/4~�;30� �EFV�XI�b< @%1�O㠮3� _RT;RQ��= D�`@���Q@  �EjP"�㥎�<�B�� <	�@��AMP��]>�a�����a�8S�q�DU�@q���"C�AB��?A��0NSls���IDI�WRK�h^�� V�WV_]�~��> �DI��q�@� /.�L_SE2�T���/��Z`��0��#�E_п�u�v�j��SW�J�j� 𲰂�	���=�c�OH�z�PPLJ�v�IR!��B� ���w�d��B"����BASh��� X ���V�����?C��Q��R7QDW��MS����AX}�8�u�LIFAE� �7�A1C�NJ� ��S��H���Cs�>�Z�C`QN"䘡U��OV� _�H9E����SUP�hb�C�� _�Ԥ���_P����[Q��Z��W����ו�Tb��XZX$ `1��Y2F�CM@�T��t@�N�p�	8�!��9A `�P.�sHE��SIZy���u��BN�pUFFI���p� �Q/4�0�<2671�!MS�W9B 8�KE�YIMAG�CTM�@A��A�Jr�>�!OCVIET���'C C�V L�t����s?� |� :D��"pST�! x�0�� 0��Ѡ��0�>��EMAIL���@���g0c`_FAUL⍢EH�CCOU��p}$T@��F<' $���eS]���;ITvBUF��qP���T  ���B�dC�t����#��SAVb$)�e�A� }���Pi�e@U��b`_ H���	OT{BH�lcPր(0�
{��AX1#�� @��_GJ�f1YN_�� Gj�D�U/0eU��M����T8��F��ِ�A!H��(@u���C_r@�@K�D����=p�R���uDSPl �uPC�IMb ��J���U����Eƀ��IP�su��D`�TH0�c���TuA�HSDI�ABSC�ts��0Vzp*} �$�#��NVW�G�#�$0� FJ�/d�jƓASC��U�ME�R��uFBCMPL��tETH�!AI��FU��DU �a�@;⠂CD�O � ����R_NOAUT.g` J��Pp2X��n4ĥPSm5C`%}5CI�.ak3|� =KH *}1Lp��Q��&�I� ��4#Q�6s��6ѡ�6P0��6���67�98�9�9�:J��8�:1J1�J1J1+J18J1�EJ1RJ1_J2mJ2T�;J2J2J2+JU28J2EJ2RJ2_J�3mJ3�:3KJ3PJ/�G8J3EJ3RJ�3_J4mB���EXT�>aLC` ��F�fF�5Q9g�5���FDR�MT��VC��C�wa}".C�REM,�FAj�OVM��eA�iT7ROV�iDTm �jMX�lIN�i���jN�IND�`!�
x<p /$DG�Ð�`opS�9�D��`R�IV)0Qbj�GEA-R�IO0�K�bu�Nj�x�.؎��p�q>j�Z_MCM>�C��d`��UR)2N ,<{1��? ��
 s?�pI�?�q�E���q0�T0lbOԁ���P� �RI�T5��UP2_ gP Ѡ#TD=  ��C����qP�J�6�$wBAC;Q T��h$9 O�)��OG���%E��3e&0IFI���e0�0����PT��caMR2ieRO vbY�vbLIq��{g���P�f��Ŗb_mAN~"F�_F�I4+�M;v`�r}DGCLF��D7GDY��LD�q>tA5[�5S�كk�S���M� T�FS� l�T P�)���|
�/$EX_)��@�)�1�� ��*�3�b�5b��G�!ieU� � p&2SWKO>��DEBUG�S���0�GRY�zU�#B�KU� O1�@ O�PO8��Π0l��ΠMS]�OO��SM]�Eq��p�Q`_E V �$�X� �TER�M2�W;�`��OR�IĀ6�X;����S#M_��$7�Y;�#���TAy�Z;� ��UPB�[� 9-��QbV$G����W$SEGźאE�LTO��$US]E0NFI�����p���`���X$UFR����q0豈�D5fh�OT1Ǵ TA_ ��C�NSTd�PA�TT!��Y�PTHJ�!B0En�K0�ART� ���������REL��&SHF�TF"�_���_SH"��M�!B0x� ��n�r��Z���OVR
#N&SHI����U�2= �AYLO$ 5I1�_�d���d�ERV�0*�} ��b ?�d��Q����A���RC
���ASYMh���WJ�apAE�����f�2�U��@d�5����D5��P#XGи!	�ORd�M�&��GR!���\��΢��^�����k�]� �E���TO�C�졳q��OP@��N z�3&1���aYO�a> RE��R�#b&O0��`�e���R]��������e$7PWRSpIM��[�sR_���VISy��r���UD�t�� ;^>�$H����__ADDR9fH$�AGa�z�s�i1R\� =_ H8�S�  ��S��C��C��CcSE�abaHSO0���` $���_aD`���PR�w�1HTT� wUTH�a ({0�OBJE1u���-$9fLEP�-=�b � *g!AKB_qT��Sk�#DBGLV5#K�RL"�HIT�B�G0LO���TEM4$��b�������SS�p�4JQUE?RY_FLA��f QWYA���c���f� PU�"B�IO0 ��4G��H��HB� �IOLN~�d�/0i�C��$S�L�� PUT_&�$���Pwp��rSLA�� e /2����ӡ��,�{IO F_AS�f��$L��U�� �#�04�#����,��HYOgN!'#�UOP�g ` l!9f@�b>$�`E&�!��P�����'�!E&�"�&؁I�P_MEMBk0T� h X IPz�v��"_#0v�����0��Oc6�1w�DS�P�' $FOCUgSBGv��0UJhf�i � 60S��JsOG�W2DIS��J7��O��$J8�97��I6!�2�77_LABQ����0��8�1APHI�p�Q�3�7D+�J7JxRA4`P�_KEYp� �KILM�ON�j&`$X�R =0cWATC�H_ �DӘ�U1EL�� �yc`B�k �GpG�VP�-ffBCTaR��fB5baLG|�l ��+h�"��LG_SIZ{Y��E�
��F
 �FFD�HI �H�H��F�HM��F�@ ���C5V
�5V
 5V�@5VM�5W�`S)@S�����@Nv1��mx �� ��R��4a�PÀU��Qk�L�S�RDAU�UEA I���R��PGH��r� BO}O~�n� C-"�2�ITGcd��)&R{EC-jSCRN�)&DI(#S��RG����cl�!#��b$�!Sa"Wkd!ܽT!#JGM�gMN3CH"FN�2�f�K�gPRG�iUF��h	��hFWD�hH]L/ySTP�jV�h�Ā�h`�hRSgyH!�{&C�Es��!#���g�yUt�g��f|@6#�bG�i4�P!O�JzZeEsM�w82v�iEX'TUI�e	IP�cw��c���c ���`�a����s��Jg���KaNO{�ANA8"貇�VAI�0z�CL����DCS_CHI��������O�L���SI)��S'��hIGN�@��C�arT����DEV�wcLL�єQ6@BU𠪔�oa@�T��$�GEM'9nDdѢ��pa@ЅC\�!��OS1��2���3��*3�����q �T0v-�絡.e�IDX���-f�L�b�STm R�PY�0���� p$E��C���  ����8� ��r L*</���Q(6����6�EN� 6�ՕKc_ s Y��P$ dKaD�� �MC�Rt =�T0CLDPm ��TRQLI`��e0x�f�FL>1��_���b�DUA��LD������ORGe0�r�� �WX�����Y���V�O�?u � 	���u�u���Si�Tx��0�0�ްS�[�RCLMCi����{�m[��ՐMI��O�v d��Q6�RQ�00�DgSTB��Y� ��{a��AX��@�� �_EXCES����)M��wA0�¹�Q����x(��_A�ʊ l����V�K|�y \*�2��7$MBLIE��?REQUIR��z��O��DEBU*��L�M{�zW�.!P��B��i���N,0�3Ѩ�{�R�RkHV�DCE��TIN3 `!�TGRSMw0p�S�N������s<�PST�  �|h�LOC9�RYI� 9�EX��A��x:�����ODAQo%�}��$@�Q΂MF�A�_���p�8C��P��SUP����FX��IGG�"~ �0��MQ���v�5@� %����m ���m ����6#DAT	A����E� 1�NP�" N�� t�MDIF)?�!��H���1!� �1"ANSW�a!ܑS�!D�)��H3Q�n$� ?�CU�@aV_ >0���LO�P"$�=ұ���L2т�����RR�2I5��  ��QA�X� d$CALII��NUG�2g�RINp<$R�SW0��K�A�BC�D_J2SqE����_J3v
p1SP�@6 ��	Pp�3��\�����J���P�O村IM��[�CSKAP��$�P�$J�Q[�Q,6%%6%,'���_AZW��h!ELx�����OCMP�����1X0RT�Q�#�c1�c@�Y�1��(t�0�*Z�$SMG�p�����ERJ�ԑIN� ACߒ�@�5�b��1�_B��542d���14X҆f>9DI~!��DH �t30���$Vlo�Y�$�a$�  ��A�<�.A�����H �$BE�Ly lH�ACCE�L?��8���0IR�C_R��&��AT<w�c�$PS �k�L͠yP D��0Gx�Q�FPATH�9�WG�3WG3&B��#�_@�2�@�AV���C;@��0_MG|a$D�D�A@[b$FW�(����3�E�3�2�HD}E�KPPABN.GROTSPEE�B���_x�,!��DEF�g��1͠$USE)_��Pz�C ����YP�0V� �YN���A{`uV�8uQM�OU�ANG�2�@O9LGC�TINC~����B�D���W���ENCS����A�2��@INk�I&Be���Z�, VE�P'b2�3_UI!<�9cLOWL3��pc x��UYfD�p��Y�� ��Ury�C$0 fMOS`�Ɛ�MO����V�PE�RCH  vcOV�$ �g9��c��\bYĀ���'�"_Ue@0��A&BuL������!epc�\jWvrfTRK�%h�AY�shчq&B��u�s���&l��Rx�MOM|���h�ﰞ �Ą�C�sYC���0D�U��BS_BCKLSH_C&B��P �f�`}S�7��RB��Q.%CLAL��b?�8�pX�t�CHKx�H��S�PRTY�����e�����_~��d_�UMl�ĉCу�ASsCLބ PLMT��_L�#��H�E ������E�H�`-��Q#p_��hPC�aB�hH��ЯEǅCw���XT�0�GCN_b(N�þ���SF�1�iV_RG�e�!��&B����CATΎSH ~�(�D�V��f�0'A�	� �@PA΄�R_Pͅ�s_y�뀎v`�`x��s����JG5��6Ф�G`OG���rTORQUQP��c�y��@�Ңb�q�@�_W �u�t�!�14��33��3�3�I;�II�I�3F��&������@VC"�00���©�1��2�8ÿ�¶�JRK�����綒 DBL_SMt�QO�Mm�_DL�1O�GRV:�3ĝ33��3�H_��Z@a��COSn˛ n�LN ���˲��ĝ0��� �� e��ʽ̃��Z���f��MY���z�TH|��.�THET0beNK23�3Xҗ3��[CB]�CB�3C��AS���e��ѝ3���]�SB�3��h�GT	S@! QC���'y�x�'����$DU�� ;w	��Q�����q9Q����$NE$T�!I�����)I7${0LсAP�y��`�k�k�LCPHn�W�1eW�S�� �������W���������{0V��V��0��UV��V��V��V��UV��V�V�H��@����7�����H��UH��H��H�H��O��O��OF	��O���O��O��O��O*��O�O��FW�}���	�����SPBA�LANCE�{�LmE��H_P�SP1��1��1��PFULC5\D\��:{1��!UTO_���ĥT1T2��22N���2, ����q^P<�-B#�qTHpO~ |�1$�INSEG�2�{aREV�{`aD3IFquC91�('o21�dpOB!d�=���w2��7P���LC�HWARR�2AB����u$MECH`��ДQ�!��AX�q�PB��&r�~2�� �
�"��1eROBƬ`CR r�%���?�MSK_�4_� P �_OPAR�1�2(47Qst1��,`*R(0)cB�(0|!I�N!�MTCO�M_C���0� � �@0 �A$N'OREc�2�l ~2o� 4�GR��%FLA!$XYZ_DA��LP;@/DEBU�2 �0lR֫0� ($mQCODS� �2�r� ��p$BUFI�NDX*P �2M{OR3� H%0 �p�0��:@�p�QB�"��1��NF�TMA9Q#C�rG.B�� � $SIMUL���0�As�A�sOBJE3�FA�DJUS�H�@AY�_I��xD�GOU�TΠ�4�p�P_FI�Q=8AT#�Y,` W�1P +�PQ+ 9�:uDjPFRI �PUMT0�RO�
`E+�>Sp�OPWO��0��,@SYSByUi� @$SOP�Q�By��ZU�[+ PR�UNn2�UPA;0D�V�"�Q�`_�@F��P�P!AB�!H��@IMKAGS�%0?�P!3IMQAdIN$��R~cRGOVRDEQ�R�@�QP�Pc�� �L_��feÂސR�Bߐ<pX�MC_SED'@�  H�Ni �M�bG��MY19�F�#@EaSL30�� x $OVS�L�SDIsPDEAXǓ�f֓Hq�bV+��eN�a
��Pp�cw�x�bw��d_SE9T�0� @�CrL�%9�RI�A3�
Vv!_��bw{qnq#@-!\�@� �4BT� �àATUS�$�TRCA�@PB�sB�TM�w�qI�Q�d4pF��s�`0� D%0!E�P�b�rr�E1"�qpQpd��qEXE�p@���a�"��tKs�Rp�&0�pUP�01�$Q `XNN�w���d����y �PG|5�� $SUB�q�%xq�q|sJMP�WAI$�Ps��L�O ��1
 �E$R�CVFAIL_C@1�PÁR%P�0�#����Ȕ� �
�R_P=L|sDBTBá��ΧPBWD��0UM��IG�Q `�,�GTNL ��b�ReQ��2���qP��@E�Ǔ��֒��DEFS}P� � L%0ĺ ��_���CƓUN!I�S�wĐe�R)���+�_L
 P�q�#@PH_PK�5�~�2RETRIE|s̛2�R���FI~�2� � $��@� 2��0DB�GLV�LOGSCIZ�C� ���U�"2|�D?�g�_T:��!eM�@C
 #EM���R��y0�8CHEC�KS�B�Po01�B�0.�0R!LbNMGKET��@�3砹PV�1� h�`A�Rp� �1)P�2>�S��@OR|sFORM3AT�L�CO�`q�d���$Z��UX�P�!r�LIG�1��  ˣSWI�m �a�q��,�G�AL?_ � $`@R��B�a��CS2D�Q�$E1��J3�DƸ� T�`PD�CK�`�!LbCO_J3����T1׿6� �˰C_Q�`� � ��PA�Y��S2u�_1|�2|�ȰJ3�ИˈŬƼ��tQTIA4��5:��6S2MOMK@�à��������y0B׀A�D��������PU��NR��C���C�������4�` I$PIN�u�41�ž� ��:q�R~ȇ��ٯ� �:�h��a�֬��ց��1�'1R\uSPEED G��0�؅�� 7浔؅�%P7�m�F�p�U��؅SAM �=G��7��؅MOV	B� e0�� ��c2 ��v��浐�� ���c2@nPsR����İ$QH���IN8�İ��?�[��6�؂A���X����G�AMM�q�4$GGET1R@�SDe�zmB
�LIBR[��y�I�7$HI�0_�5a@c2E`@#A@ 1LW^U�@	�1a¬&o�ʱC�=�n S`�p �I_��pPmDòv� ñ'����mD��	ȳ� �$�� �1��0IzpR� D`T#|"c���~ LE^1�41�qwa�?�|�M�SWFL�MȰSCRk�7�0��Ѻpv���Z 0�P�@�9@���2�cS_SAVE_Dkd%]�NOe�C�q^�f�  ��uϟ�}ɕQ��}��Ѐ}*m+��9��ժ(��D �@���������b3 1�RA�Mam�7
5�#���^���Mtա 7� �YL��
A
'�VAS	BtRna`7 GP�B
Bl3
A%`�$GSB1W? �2�2c�Ȭ3oBB1M&@�;CL �8���G�b�1v���9M!Lr� �N�X0�d$W @�ej@b �� @=�BD�BK�B �-�> �P����ycJİX �OL�ñZ�E����uԣ ��OM�R/d/v/�/ �/��A�jM`��e�_��� |��H  ��jV��yV��yP�ʗW�V��E���
�MS������NTP=���PMpQU�� �� 8TpQCOU�,�QTHQ�HO�Y2`HYSa�ES���aUE `"#�O.���   �P�0��rUN�p�3��O$�J0� P�p^e��x����OGRA�q�k22�O�d^eITxm�aB`INFOI1����k�ak2��O�I�b� (!SLEQ(��a��`�foayS� ��� 4Tp�ENABLBbpPTION|s����Yw���1sGCF��O�c$J�ñfb���R�x!�]ot�bS�_EDŀJ0� ��N��@K�᪃E�S NU�w�xAUT<,!�uCOPY����(�v�8 MN��^�PRUT�� ��N�pOU��$G�cbn��aRGAD5JI1�2�X_B0ݒC$ ����@��W���P�����@㊀��E�X�YCLB��RG�NS6u�N0�LG�O�A�NYQ_FREQZ�W���+�p�\cLAm"�������uCRE  c� �IF�ѝcNA���%i�_GmSTA�TUQPmMAIL�� 1��yd�����!��ELEM��� �7 DxFEASIGq2��v��q!�er$�  I�`�"�`�ae�|I�ABUq��E�`D�V֑a�BCAS��b� [�Ub��r % $y���RMS_TRC�ñj ���Ca��ϑ��,r����C�YP	 � 2� g�DU�� ���Ԣ�0-�1��1����qDOU�ceNLrs��PR30;p�r�GRID�aUsBA�RS(�TYHs��O�TO�I1��P`_"��!ƀ��l�O�@7t�� � �`�@P�OR�cճ��ֲSReV��)���DI. T���!��+��+�U4)�5)�6)�7)�I8��aF��:q�M`?$VALU|�%��ޡ��7t�� !Cu'!�a���� (FgpAN#��R�p|0� 1TOTAL��,[��PW�It�&�REGEN$�9��S�X��sc0��Q���PT1R��Z�$�_S ��9дsV���t���rb�E��x�a�"^b�p��7V_H��DA�C�Ў��S_Y4!�B<�S��AR�@2� >f�IG_SEc��d�˕_b`��C_����w��?r��%�b�H�SLG#�I1��p@"=���4��S�2̔DE�U!Tf.p��TE�@����# !a����Jv�,"��IL_MK��z�н@TQ�P�a��T��2VF�CT�P���^�Mu�V1t�VU1��2��2��3��3��4��4����������1�"IN	VIB@N�; �!�B2>2J3>3
J4>4JI05����"���p�MC�_F`3 � LP!!�r�M= I���M� [PR��� KEEP_HNADD�!f�	C�A��!����"O�Q I����"���?�"REM9@!�ϲ^uzU���e!HPWD  �SBMSK"G�a	!B2B�
#?COLLAB�!@��2�����o��`�IT��A`��D�� ,pFLI@��O$SYN� ;,M�@�C>��%�UP_D�LYI1�MbDEL�Am ј�Y�PAD��A�qQSKIPNE5� ��``On@cNT�1� P_`` �b�'�`�B]0�'���) 3��)��)O��*\��*@i��*v��*���*9O�J2R‎��?sEX��T%�|1�{2�ܐ�|1�a���wRDC!F� ��pER�sR�PM�'R^�p�:b�2�RGE�p82��3d�FLG�Q�J��t�SPC�c�U�M_|0��2TH2�NP�F@o0 1��  �x��p11��� l[P�E-Ds#ATWo�[�w �B�`�d�A�p3�BfcBAHnP�B��_D2gB�mOO�O�O�O�O�G3gB��O�O_ _2_D_�G4gB�g_y_�_P�_�_�_�G5gB��_@�_oo,o>o�G6gB�aoso�o�o�o�o�G7gB��o�o&8�G8gB�[m�����ES����\@ǡ`CN�@�_@ZwE��^� @�o��m�IO�ፉI����j�POWE!� W�: �18���0� �5%Ȃ$DSB;���֒ ��h CL@�Г!RS2;32s�� ��0�uy.��ICEU{�暐PEV@��PARsIT�њ�OPB ���FLOW�TR`2�҆]���CUN�=M�UXTA����INTERFAC�3�fU���CH�� t� � ˠ�E�A$����OM$��A�0נI����/�A�TN����Tо ��ߓ��EFA�� �"!�Ґ�� Hu!��� O�� &�*�� �����  2� �S�0~�`�	� �$3@B}%:B�Ŏ��_�DSP��JOG���V�h�_P�!s�OANq0%�0���K���_MIR���w�MT7��AP)�w�>@"���;AS������;A{PG7�BRKH����G �µ! ^���i��P��Ҏ���BS�OC��wN���1�6�SVGDE_�OP%�FSPD_�OVR�u �DLвӣOR޷�pN��b߶F_�����OV��CSF�<��
�F0Ƽ���UFRAF�TOd�LCHk"%�#OVϴ ��W[ ����8�Ң�͠;� ; @ BTIN����_$OFS��CK��WD���������r,���TR��T��_FD� �MB_)C �B��B��0��(�.Ѻ�SVe�Ґ琄�}#�G)�<�AM��B_��jթ߃_M@�~��ቂ��T�$CA����De����HBK�����I�O��թ���PPA��������Տթ�~��DVC_DB�� ?����A��,�X� b��X�3`���3�0�����ϱU󳠈�CAB�0��ˠ��c�� �Ow�UX��SUOBCPU�ˠS�0 �0�R����!�A�R��ł�!$HW_C@g@A��!��F��!�p�� � �$U r�|l�e�ATTRI���y�ˠCYC����C9A���FLT ��`������ALP׫�CHK�_SCT6��F_e�F_o���Ɓ�FS�J�j�CH�A�1��9I�s�8RSD_!聂��恩��_Tg�7�� �i�E)M,��0Mf�T&� �@�&�#�DIA�G��RAILACN���M�0�"��1`���L��{�PRB�MS   �pC4�z&�	��FUNC�"���RIN�0 "$0�7h�� S_��(@��`�0��`A��GCBL� u�A����DAp�a���LDܐð���d��j��TI�%��@�$CE_gRIAA��AF��P=�>#��D%T2b� C��a�;�OIp��DF_Lc�X�葶@�LML�FA��H�RDYO���RG��HZ 7����%MULSE� �����.k$JۺJ�����FAN_ALMsLV�1WRN5HARDr��Fk�2$SHADOW |�A���O2s�0N�r��J�_}���AU- R�+�TO_SBR ���3���:e�6�?�3_MPINF@{�8�4��3REG�N1DG�6CV��s
��FLW��m�DAL_N�:�����q��	����a�U��$�$Y_Bґ� u�_�z��� �/�EGe���ð�A#AR������2�Gܷ<�AXE��RO�B��RED��WRd��c�_�M��SY`���Ae�VSWWRI���FE�STՀ����d��Eg�)��D-�	{2��BUP��\V��]D��OTO�1)���ARY���R����6�נFIE���$�LINK�!GTH��R�T_RS��8�E��QXYZ��Z�5�VOFF���R��R�X�OB��,`8d����9cFI��Rg��􃻴,��_J$�F�貿S��q0kTu[6��1�w �a�"�b�CԀ+�DU�¤F7.�TUR0X#�eġQ�2X$P�ЩgFL��Pd���@p�UXZ8����� 1�)�KʠM��F9���ӓORQ���f&ZW30�B�OPd��,��t����A�tOV	E�qeBM���q^C�u dC�ujB�v�wL�wg��tAN=�Q�qD! fA�q��=�}��q�u�q����dC��"���ERϡj	�E��T�ńAs�@�UeX�0�W����AX��F� ���N�R��+��! +�� *�`*��`*��` *�Rp*�xp*�1�p*� � '�� 7�� G�� W� � g�� w�� ��� ��� ��đ��DEBU=�$8D3�h���RAB������sV��<� 
��i�fA ��-񷧴������a ���a���a��Rq��xq�J$�`D"�R9cLAB�Ob�u9�F�GROh��b=<��B_� ��AT�I`�0`����u8���1��ANDfp��@�����U���1ٷ �р�0�Q������PN�T$0M�SERV9E�y@� $%`dmAu�!9�PO�� [0ЍP@�o@*�c�x@�  $]�TRQ�2
\��Bf��j�D"2�{�" � ?_ � l"T�Nc6ERRub�I��qVO`Z���TOQY��V�L�@)�1R�Ƅ G;�%�Q�2 [�T0e�G� ,7�ř��]��RA#� 2� �d@����r� �Y@$�p�t ���OC�f�� � ��COUNT�UQ�FZN_CFGe�� 4B�F��Tf4;�~�\� �
��y��uC� ���M: �"fA��U��q: ��FA1 d�?&�X��@=����eB�A<�����AP��o@HEL�@��� 5��`B_BAS�3RSSRF �CSg�!��1
ש�2��3���4��5��6��7r��8
ל�ROO��йP�PNLdA�cAqBH�� ��ACK���INn�T��GB$Upq0� +\�_PU��,@0��OUJ�PHH����, u��TPF?WD_KAR��@&��REGĨ P�P�n]QUEJRO�p�`2r>0o1I0������P����6�QSEMг�O��� A�ST�Yk�SO: �4DI�w�E���r!_T}M7CMANRQ���PEND�t$K�EYSWITCH����� HE�`BoEATMW3PE�@CLE��]|� U���F>��S�DO_�HOMB O>�_�EF��PR>a9B�ABP�x�CO�!��#�O�V_M�b[0# IOcCM�d'eQ�v��HKxA� D�Q$G��Ue2M�����cFORCCWcAR�"̀��OM�@ � @r�:#�0UUHSP�@1&2&&E3&&4�A��s�O���L"�,�HUNLiO��c4j$EDt1�  �SNPXw_AS��� 0+@� @��W1$SIZ��1$VA���M_ULTIPL��#�! A!� � �$��� NS`�BS��ӂAC���&FRI	F�n�S��)R� {NF�ODBU$P����%B3=9G�r��Sܪ�y@� x��SI���TE3s�r�cSG%L�1T�R$p&�П3xa�P�0STMT1q2�3P�@5VBW�p�4�SHOW�5��SmV��_G��� Rp�$PCi�oз��F�B�PHSP' A�v�Eo@VD�0vC��� ���A00 ޴RB% ZG/ ZG9 ZGTC ZG5XI6XI7XIU8XI9XIAXIBXI@ ZG3�[F8PZGFXH���XdI1qI1~I1��I1�I1�I1�I1��I1�I1�I1�I1��I1 Y1Y1Y2�WI2dI2qI2~I2�I2�I�`�X�IQp�X��I2�I2�I2�I2
 Y2Y2Y�p�hdIU3qI3~I3�I3�IU3�I3�I3�I3�IU3�I3�I3�I3 YU3Y3Y4WI4dIU4qI4~I4�I4�IU4�I4�I4�I4�IU4�I4�I4�I4 YU4Y4Y5�y5dIU5qI5~I5�I5�IU5�I5�I5�I5�IU5�I5�I5�I5 YU5Y5Y6�y6dIU6qI6~I6�I6�IU6�I6�I6�I6�IU6�I6�I6�I6 YU6Y6Y7�y7dIU7qI7~I7�I7�IU7�I7�I7�I7�IU7�I7�I7�I7 Yu7Y7T��0�P� Uc�� �l�נ��
>A820��j���RCM2����MT�R��|���Q_��R-��ń�����[�YSL�1�� � �%^2��-4�'�4��-Y�BVALAU�Ձ���)���FJ��ID_L���HIr��I��LE_������$OE�SA~b�� h 7�VE_BLCK�¡1'�D_CPU 7ɩ 7ɝ �����E����R � � PW��>�E ��LA�1Saѝî����RUN_FLG �Ŝ������ �����Ą����H���Ч��}�TBC2��� � _ B��� b�r� W?�eTDC����X��3f�S�CTHe�����R>�~k�ESERVEX��e��3�2 �d���� �X -$��LENX��e����RA��3�LOWI_7�d�1��Ҵ2 �MO/�s%S80t�I���"�ޱH����]�DyEm�41LACE��2�CCr#"�_M�A� l��|��TCV����|�T�������0Bk�)A�|�)AJ$��%EM7���J��B@Rk�X�|���2p `�0:@q�j�x JK��VKX�����ы�J0����JJ��JJ��AAL���������4��5�Ӵ NA1�� ����LF�a_�1� H! �CF�"�� `�GROUP���1�AN6�C�#~\ REQUIR�Ҏ4EBU�#��8�$Tm�2���|�ё %�� \�A�PPR� CA�
�$OPEN�CLOS<�Sv��	k�
��&� �<�M�hЫ���v"/_MG�9CD@�C ���DBRKBNOL�DB�0RTMO_�7ӈr3J��P ��������������6��1�@ �	�$��� � ���'��-#PATH)'B!8#B!��>#� � �@�1S�CA���8INF��UCL�]1� C2@UM�(Y"��#�"������*���*��� PA�YLOA�J2L�ڠR_AN`�3L���9
1�)1CR_�F2LSHi2D4L�O4�!H7�#V7�#ACRL_�%�0�'��$��H���$H�C�2FLEX�:�J#�� P�4��F߭߿���0��� :����|�HG_D�����|���'�F1 _A�E�G6�H�Z�l�~����BE�������� ����*��X�T,�C� ���@�XK�]�o�^Av�	T&g�QX>�?��4T X���eoX�������� ����������	-	:"J@� �/�M0_q~�۠AT�F��6�ELHP���s�Jڗ � JEoCTR�!�ATN���v|HAND_VB�q�1��$� $:`�F2Cx���SW�Ms��� $$M,00�_Y�n i��P\����A��� 3����<AM��_AmA|��NP�_UDmD|P\ G���E�STaM�nM�NDY��� C���� 0��>7_A>7Y1�'��d�@i`�P���@����"��J$�� O�4D'"��J�<��ASYMl%A�	� l&��@�-Y1�/_�}8� �$��� � �/�/�/�/3J	<��:;�1�:9�D_VI��x���V_UCNI�ӝ��cF1J�� ��䕶�Y<��p5Ǵ� y=6��9��?�?>�wc��4�3  �$�� ASS  ����s�=�=� �h�VERSIO�Np�~��=
��IRTU<�q����AAVM_WR�K 2 ��� 0  G�5z�������.� �	8�)�L�=����:�w�^�|�(ܛݧ�7ѭ�����|����BSPOS�� 1��� <��A�S�e�w� ������������ �+�=�O�a�s����� ����������' 9K]o���� ����#5G Yk}����� ��//1/C/U/�>��AXLMT��X#��%�  dj$I�Ns/�!i$PRE_EXE�(� �&)0�q�������LAR�MRECOV ��ɥ"
�LMDG� ����[/LM_IF �� �!X/c?u?�?�?�:Q?��?�?�? OM, 
0�8O�4�cOuO�O��O�NGTOL � ���A   ��O�K��PP)�O ; ?6_,_>_P_{� $BR_�_ w�o_�_�_�_�_�_o@�_'oo7o]o�!��O �o�o�o�o�o�o�o�+=Oa�PP�LICAT��?��� �%@�Handling�Tool �u �
V8.30P/�33�@lt��?
88340�slu

F0�q��z=�
2026��tlu��_�7DC3�p�J  �sNone�lx� FRA������B��TIV�%�s�#~��UTOMOD� �E�)P_CHGAPON������Ҁ�OUPLED 1��� ��"��4�uz_CUREQ7 1��  � >�>�*ސ�4��!���x�~� ��u��Hm����HTTHKY�� ��w���7����%�C� I�[�m��������ǯ ٯ3����!�?�E�W� i�{�������ÿտ/� ����;�A�S�e�w� �ϛϭϿ���+���� �7�=�O�a�s߅ߗ� �߻���'�����3� 9�K�]�o����� ��#������/�5�G� Y�k�}��������� ����+1CUg y������ 	'-?Qcu� ���/��/#/ )/;/M/_/q/�/�/�/ �/?�/�/??%?7?�I?[?m??��P�TO��@����DO_CL�EAN܏��CNMw  �K >��aOsO�O�O�OD�DS�PDRYRO̅H	I��=M@NO_'_9_ K_]_o_�_�_�_�_�_8�_�_J�MAX�p�4�1���aX�4"��|"���PLUGG����7���PRC�@B�;@?K_�_ebOxjb�O��SEGFӀK�o�g�a;OMO'�9K]�o�aLAP �O~Ǔ����� ��/�A�S�e�w���>΃TOTAL-fVi�΃USENU�`��� ��䏺�P�RGDISPMMC�`e{qC�aa@@}r���O�@f�e��_�STRING 1�	ˋ
�M�ĀS��
`�_I�TEM1j�  n ����������Ο��� ��(�:�L�^�p����������ʯܯI�/O SIGNA�Ld�Tryout Modek��Inp�Sim�ulatedo��Out.�OV�ERR�@ = 1�00n�In c�ycl"�o�Prog Abor8��o��Statu�sm�	Heart�beati�MH� Faul����Aler���ݿ�π�%�7�I�[�m�� �3f��1x����� ������*�<�N�`� r߄ߖߨߺ�������8���WOR�`f� L���&�t����� ��������(�:�L��^�p�����������POd�����d��� %7I[m�� �����!3pEWi��DEV�� ������/ /'/9/K/]/o/�/�/��/�/�/�/�/�/?PALT��81d�? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnOp�O�O�O&?GRI` f��AP?�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHo�OR�̀a�OZo�o�o �o�o�o&8J \n������<�noPREG<>%� �o�L�^�p������� ��ʏ܏� ��$�6��H�Z�l�~�����$�ARG_L�D ?�	���ӑ��  	�$�	[�]�����ƐSBN�_CONFIG S
ӛ&�%� ��CII_SAVE  �E�<�Ɛ�TCELLSET�UP Ӛ%  OME_IO���%MOV_H8������REP�l����UTOBACK�t�0�FRA;:\� ����_�'`���=�{� J� 	� �����ͿĿֿ�6����	�1�C�U�g� yϋ��Ϸ������� ��ߜ�5�G�Y�k�}� �ߡ�,���������� ��C�U�g�y���\��a�  )�_��_\ATBCKC�TL.TMP DATE.D;<��	�p�-�?��INI;0�p�8��MESSAGT�^�_�ېi�ODE_D��W�8��H���O����PA�US��!�ӛ ((O֒��
�� *N<r`�� �����"��~��TSK  ��x=�C�	�UPDT���\�d���XWZD_ENB\�4���STA[�ӑ�őX�IS&�UNT 2�ӕ`� � 	�S��c2��V0�D�[*� Q����  %�`'$h�
/L/�^. "YK��ާJ'"��b}�2c/�/_/�/��/�MET�`2��P�/?�/<?�)S�CRDCFG 1�C`��\�\�1?�?�?�?�?�?�?6��QX��??O QOcOuO�O�O O�O$O �O�O__)_;_�O�O���GR����zS���NA��қ	��wV_EDZ�1ze9�9 �%-��EDT-h_ʪ�_o&�`/A���-��_
�	������_�o/  ���e2�oɫ ko�o�6k�o!hozo�o�c3Y�o��o �n��4F�j�c4%��r���nN���  ����6��c5�a� >����n���̏ޏt���c6��-�
�Q��n��Q�����@�Ο�c7 ����֯��n���d�v�����c8U��_����0
 }~��0�B�ؿf��c9!ϑ�nϵ� }Jϵ���Ϥ�2��aCR�oį9�K��� ������n���zP�P?NO_DEL�_xR�GE_UNUSE��_vTIGALLO�W 1�Y~�(�*SYSTE�M* 3	$SERV_GR�R 69�n��REGB�$d� <9�NUMg��z��PMU�� 5�LAY�  <�PMPAL[��COYC10������<����ULSU��{�����D�L�N�B�OXORIk�CU�R_;�z�PMC�NV��;�10|���T4DLI�4�V���ߨ�� '9K]oR�zP�LAL_OUT �Dcc�QWD_�ABOR��	��I�TR_RTN��<�Y� NONS8�� �CE_RIWA_I��<�F_1��B =�[_PARAMG�P 1��w`_����CWp  .� � U� � � � U� � � � �� � �  DF5`D$3!g-�<$��H$�T$� DUX � X "� �B�D1� 9X @�� 6?� <HE��O�NFIy���!G_�P��1�  �e�U??0?B?T?f?�x?�?�!KPAUS�X�1�UR , Z��?�?�?�?�?OO OTO>OxObO�O�O�O��O�O�O_�2O_�ey�PCOLL/ECT__�Y5auGWEN��I�"cRn QNDEOS�W���1234?567890�W��S�u�_�Vy
 H�y)�_#oS��_o hoT�AoSo�owo�o�o �o�o�o�o<+ �Oas���� ����\�'�9�K����o��VQ�2W[� � t�VIO �YcQyH&�8��J�\��TR�2؍(��
��j�� � ����%�_M+OR҂!� + �'� 	 �5�#��Y�G�}�k����Ӂ"��2?�!�!3 ҡR�Kڤ��$R_�#*_	���C4 c AS yC  x�{A3!z  BC!��PB/!�PC  �@*����:Wd�
�IPS$����T��FPROG %�*6߼�8���I����&RҴK�EY_TBL  �)VR� �	
��� !"�#$%&'()*�+,-./�W:;�<=>?@ABC���GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾���������͓��������������������������������������������������?�������1���LCKۼ3���S�TA�д_AUT���O(��U�IN�DtTD�FQR_T1_�Q�T2��7$��6��XC� 2�����P8
SONY? XC-56�������@����u� ��А�HR5��cT0�B�y7T�f�Affr������� ������� 5�G�"�k�}�X��������������ǼT{RL��LETEG���T_SCRE�EN �*�kcsc:U$MMENU 1&�)?  <�� �y��Ã� =&sJ\�� �����'/�/ ]/4/F/l/�/|/�/�/ �/�/?�/�/ ?Y?0? B?�?f?x?�?�?�?�? O�?�?COO,OyOPO bO�O�O�O�O�O�O�O -___<_u_L_^_�_ �_�_�_�_�_�_)o o o_o6oHo�olo~o�o �o�o�o�o�oI  2X�hz���� _MANUAL�߆��DB��L+�DBG_ERRL��s'�� ��\�n����NUMWLIMK�d ��p�DBPXWOR/K 1(�I�ޏ�����&�ŽDBT;B_@ )���ꌑ��qDB_�AWAY�_�GwCP  �=�װ�~�_AL��D�z���Y��M � �_)� [1*�����
͏����6�@�_MM{�ISAЉ�@B��P�ONTIMJM� ��p�ƙ
��ۓMOTNEND�߿ڔRECORDw 10}� �>�?�G�O����?� ��2�D�V�h���p��� ���*�߿�Ϛ��� 9Ϩ�]�̿�ϓϥϷ� R���J���n�#�5�G� Y���}��ϡ������ ����j���C��g� y������0���T� 	��-�?���c���\� ���������P��� ��;��_q���� �(�L%� 4[����� ^t�l!/�E/W/ i/{//�//�/2/�/��/??�/z�TOL�ERENC��B��В��L���CS�S_CNSTCYw 116�  ?Β�?�?�?�?�?�? �?OO&O8OJO`OnO��O�O�O�O�O�Oc4D�EVICE 126� b�*_?_Q_ c_u_�_�_�_�_�_�_�?�d3HNDGD �36�Cz�^L/S 24]�__o qo�o�o�o�o�o�_e2�PARAM 5��B��t�dc4SL?AVE 66�e_CFG 7���gdMC:\�e0L%04d.CSV�o��c|�r�"�A �sCH�p&a�&��n��w��f��r����ÀJ�P�>��\_CRC_OUT 8U�����oEpSGN �9U�Ƣ��\��16-OCT�-22 14:2y1�p�02���4��9V UB�u1�݁�nހ��o���Im��P��uG��@uVERSION ���V3.5.1�1E�EFLOGI�C 1:ݫ 	6��|�C���^��PROG_ENBp����͢��ULS{�� ��^�_ACC�LIM|���Xs��WRSTJ�N[���ţ�^�MO�¡Zr,�INIT� ;ݪs5� �*�OPT$p ?	�i�B�
 	Rg575�c��74��56��7��50��R��Ƣ2��6��X�y�TO  ���?�Y�]VP�DEX�d����@W�PATH ;A��A\E������7;IAG_GR�P 2@�k,��"	 E�  �F?h Fx wE?`�D��û ��V1"�ü��T0K��9�Cf�py�pY��dC�pq�B��i�ùmp�4m5 7890?123456��;�����  A��ffA�=qA���pхA��H�Aĩp�������A��Mk����@��tp�p��W0Ae�T0T0�pB4ü� Qô���
���(��A�A�
�=A�L���A���
A�Q�Au��������e������e� Pe�:�د{A�d������dѩp������Au���������r���ߖߨߺ�@�EG��A@�p:�RA5�d�/��)��#P�d�l������"�4�|F�@�Pz�AJ���c�?��9p�A3�\)A,��A&����0���������@�cP�]��AUW�P�J��C���<d�4�-d�%G��(�:�L�^�@��� $HZ��.| ����bt�  2Vh�xm������[���s�����=�
==�G���>�Ĝ��7����8��b�7�7�%�@ʏ�\"&�p�.%��@f�Ah�p9 A���<i��<xn;�=R�=s���=x<�=�~Z��;��%<'��'�~ �?+���C�  <(��U� 4"����&����%ùf��@?Œ?�?@? R?g��$^?�?"?�?�?�?�?�?�?)7L�?S�FB$�/d"Eͽ�>OG��A�Ԭq��sD�L4�x�CA��Gb�tφ���-_7_�C��_����/_�NED  E��  Eh� D�[PbRD_¿�_�86��_�_
z{_�_�w_o�K:o@bù�DP�O=�V��D@66�d��6`���A�U!o�o
o�o��o�o�o�oĿDIC�T_CONFIG; ��Yt؃�eg��ԱSTBF_TTS��
ęVs3���
�iv�[�MAU���Y�M_SW_CF*pB��s�!�OCVIEWf}pC�}����_ �!�3�E�W�i�;�� ������ȏڏ�{�� "�4�F�X�j������� ��ğ֟������0� B�T�f�x�������� ү������,�>�P� b�t��������ο� �ϓ�(�:�L�^�p�,���|RC�sDJ�r!ϐκ��������7�&�[�otSBL_�FAULT E����xu�GPMSK�_w��pTDIAG� F.y�q�I�UD1: 67�89012345��;x�MP�o!�3�E� W�i�{��������������/�A��X W!�J�"
��v�TRECP����
 �����M�(: L^p����� �� $6]�o��l��UMP_OP�TION_p�ގT�R�r`s���PM�E^u�Y_TEM�P  È�33B�pp �A  ��UNI�pau!�vY�N_BRK G��y��EMGDI_STA%�1!�rL �NCS#1H�{ @�K��9�/_}dd �/??+?=?O?a?s? �?�?�?�?�?�?�?O O'O9OKO]OoO��O �O�O�O�I�!�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXo�JO�o�o�o �o�O�o�o+= Oas����� ����'�9�K�]� wo���������oۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�o�]����� ��ɏ�����	��-� ?�Q�c�u��������� Ͽ����)�;�M� g�y��ϕϧ�]�ӯ�� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�_�q�{�� ������������� /�A�S�e�w������� ��������+= Oi�s������ ��'9K] o������� �/#/5/G/ak/}/ �/�/��/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OY/KOuO�O�O�/�/ �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oQOcOmo o�o�o�O�o�o�o�o !3EWi{� �������� /��o[oe�w������o ��я�����+�=� O�a�s���������͟ ߟ���'�9�S�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�K�9�g�yϋϥ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�C�U� _�q��9�Ϲ����� ����%�7�I�[�m� ��������������� !;�M�Wi{� ������ /ASew��� ����//+/E O/a/s/�/��/�/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�? �?O#O=/GOYOkO}O �/�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo5O 'oQocouo�O�O�o�o �o�o�o);M _q������ ���-o?oI�[�m� ��o����Ǐُ��� �!�3�E�W�i�{��� ����ß՟������ 7�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���/�9�K�]� oω��ϥϷ������� ���#�5�G�Y�k�}� �ߡ߳���������� '��C�U�g��w�� ����������	��-� ?�Q�c�u��������� �������1�;M _������ �%7I[m ������� )3/E/W/i/��/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�? �?�?�?�?O!/+O=O OOaO{/�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_O#o5oGoYosOeo �o�o�o�o�o�o�o 1CUgy�� �����o�-� ?�Q�ko}o�������� Ϗ����)�;�M� _�q���������˟ݟ �	��%�7�I�[�u� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ�a��� /�A�S�m�wωϛϭ� ����������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�e� o����������� ���#�5�G�Y�k�}� ��������������� 1C]�Sy�� �����	- ?Qcu��������� �$EN�ETMODE 1�I^� W   �(/:+
 RROR_PROG %*�%}/�)X%TAB_LE  +h��/�/�/�'X"SEV�_NUM &"  �!!0X!�_AUTO_EN�B  D%#U$_;NO21 J+9!}2  *�u0��u0�u0�u0(0+�t0�?�?�?N4HIS�3
 G;_ALMw 1K+ �u< +�?/OAO SOeOwO�O�?_2T0  +s1:"�J�
 TCP_VER� !*!u/�O$�EXTLOG_R�EQ�6�E9 SSsIZ)_TSTKFY�c5�RTOL�  
Dz�2��A T_BWD�@�P<6�Q8W_DIn�Q L^G4�8$
?"�VSTEP��_�_
 �POP_D�Oh_!FDR_G�RP 1M)B1d� 	�Ofo: W`�������g�lpw�q�ŗ��I ����fWc�o�m�o�o �o�o(L7I��m��zA�PK�A"��>�Β�� 
 E�� 	�q�@(�C��<��'�`�K�C`}dC���N��B�{���F�@UUT��UTF�Ϗj��s���s�OHcEP]���O��#M��^*�KA����?�p�F��:6:N{�r�9-�z����  �$7@��v�
�������-��+FEATURE N^��P>!Ha�ndlingTo�ol � mpB�oEngli�sh Dicti�onary�
�PR4D S�tڐard�  �ox, An�alog I/O~�  ct\b+��gle Shif�t�  !*�ut�o Softwa�re Update  fd -c��matic Ba�ckup�IF �O��ground Editސ��g R6C_amera3�F7��Part��nrR�ndIm���ps�hi��ommon� calib U䗠�n����Mon�itor�Cal�M�tr�Rel�iabL��RIN�TData ?Acquis�Z��ϠC�iagnos���0�<�almC�o�cument Viewe�\���C��ual Chec�k Safety���  - B�En�hanced U�s��Fr���8 �R5�xt. D�IO �fin� �(�@ϲend��E�rr�Lm� D �p^���s	�EN��r.�հ �P�r�dsFCTN_ Menu��v8����m�FTP I�n'�facN�=�G���p Mask �Exc��gǱis�p��HT^�Pro�xy Sv��  �VLOAאigh�-Spe��Ski^ݤ ef.>�Hf�~ٰmmunic���ons�
!
���urE�'�7�rt� F4�a�connect 2;��Incr`�str�u���� Sp�KAREL Cmod. L��ua���OAD*�=�Runw-TiưEnv�� �D;�(�el +���s��S/W�.�{�Licen�se����
����o�gBook(Sy�stem)蔭�J�MACROs�,��/Offse�S�Z�MHٰp��� wj73ΰMMR���l�35.f��e�chStop��t��R� ize*�M�i��O� 2�7�xp��0����miz���odM�witch�����a�.�� v����Optm��4q9���fil���ORD��0�g�� �8496�ulti�-T������C�PCM fun�,��.sv�o�O���� �^�5�R�egi��r��	�!�2�ri��F�  �H59k�1�Num� Sel*�  7�4 H��İ Ad�ju���adiṇ�O� ,[���tatub��\У��������RDM Ro�bot��scov�e� �d emt(�ٱn� SW��>Servoٰs��ꒄ�SNPX �b��1��g P�L�ibr���1��ڐ 9� ɰ.�30g o��tE�s�sag� f�E�@ e����"g��/I_�
�I�TMILIB���� ?P Firmn��8�^�F�Acc����<0���TPTX����510.� eln����������H5�73�rquM�i�mula��� 2n�Touz�Paxъ�1� T��6���&��ev.��I?USB po�����iP�a�� 0\�sy nexce�pt��3 <� \h�51 ����oduV#��9��Q��VN�k"6PCVL�{&�^}$SP C�SUI�d���+X�C��auҠWeb' Pl���t? �# S��\"	2��������S�&ު�V?8Gr{idplay��`&� ��8�-iRb"�.� @ � R-2�000iC/16�5¦ d+�+�la�rm Cause�/1 ed�<0:�A�scii����Lo�ad��V4�3Upl8�0�_CycL�c��m�ori����FR�A[�am�) td=t��NRTLi�3�Onݐe Hel�ݨ 542*�PC�`ρ�4�`�]�1t�rߵ48��ROS/ Ethv�t[��n�10\ҠiR}$�2D PkߵDEaR>1�E����of�AX��ΰ�FIm��F���� z��64MB DRAMު�@:�9R�FROA[�Celal3� ����shrQ�
��Zc���ÍUk�p�� pide�WteyL�s��|0\z��!CtdѰ�.��@"E7mai��li���B+�\�� R0�qZ$�GigE�N�4OL�@Sup"��b�W38oa�~�cro���� ��4��QM��Fauest�A>�j�� �miH9.dVirt`��W��0{&ImM��+T���}$Ko�l �Bui��n�յ'A�PL�&��MyV6� �"�0�*CGP�l����{RG�'p�{SKBUW�RQ�)K�&cm\:��z��fX�)�O�võ(TA�&spoҠ-�B�&��
 �I�\E P�+�CB�'fg-��&"k  �E��sv�b���vv�3��S_k��TlO;-�EH�f6.
��E�vfx_z�)�V��tr>�)�hZ%.�F�& � ��r���*�G�&���њr�����H��РJzCTIA2c�pw4�LN�1�Mr�" #[��g�""�M�-�P2�~�T�@����vxui$�-�S�&�S�&�*z4�W��2.pc�)wVGF��fxwʪ�VP2AU \fx���N�if�u���w"in��VPB����)��s�D��*��a<s�F�5 M״�s�I��c;�{&Traİ���U,p  ��<���2��RDp	�N���HY���p��-���H���Øp)����� �ϭ�����ħ���rд�<���í4+����'9L���ӎ���y�9ӫ�c<3�U��B�O�q��u��kߍӍS�y*�ߩ�\Yy<����k�W����τ�Yx����:��	������<�5�o�e/�Q�ψ�,�K�m���g��^~����u�2��A���������F��<����y�)����|����1�m�.y�+�M��8G��i�7n��c���1籖 ����yW�����7�{�����6�Z�������uk��[�|��!��?�ϔ��9iB\����_�#�{�x@.��wrst���B�� H68��@�H)T@J�EENsDI?��tql[}
_�w�P��TQ (��I)# "���PA���8T�/��85/A#bs;/�C/U/�,q �/B�Gp�/�#��/�"�36�5�R ?!2e'pai?5!:/Y48W���%INTo?e?�_.q�?4)��?�2p�a2g�?�F O��?A�ad6?��t <ZUD2gunOOqCG533R?�D�0u�O�/�Mcm���OO�LNT�?��P_�Ĕ�`0_QR7�L_�Cfi._pH?_,_f'R50�_�SAF-F�_�7�w.vo��_�_8�/�dM Cbo��̜o�bvrEo��pa�a�oaD�@�osF-AS-sS�p'Isq(�PCesXPL�O�tlo_�ut\a��Oh%afvh%- B��/����C�$��srp�?@_�?`Dw�}�bA�����h�`௏]T�ˏ�sgc�h�os�t��CG\�s;��us�?���S9g�/�G J�����GDǟi$"�o�g3diʏ!�fd����?h%J64S��Tut�o�O�?s����F�_ ����E�0���D`!�)�NO4E�O�i$3II���iwjOl�`ž��>�?*�lb
��V��vjr/��
����7��ϥ�_�?zG7\2O�EG��Ϲ?���01� ޯ��_d�oi�A8��c�50�>�x����"Lo�h%����dj9�﴿ƿؿ��c� up9�C� j�9{�E��L��Ek,B串����oS_e_��&/��O}�j94JϬ�duZ��U���=d;�����8���r7�Dhu���;]m T��������2f�a���M�`���P�-4r V���O" #S�dw�c�P�in�`�ḁ?& HTuReLf���
�?hc��g�r"��q.JG"�erM/��/ �/�LRA^��uH71��/�tCK�/<eTX�P/?i�k1/m5k.�f��riR�eH1G�/�/ cr�NNHGRf?L�iY�d7�hOuX��H\mO ��oρ�;H��DD@�O ��*�<�:I�?�?��dϜR�_ hd�gh�gOO�_���gmh�_h�m��XO�o|O�O �o�O\/�o0�f�gm�o`��`e۠;iov��yt��"��u�R60���#tm�o_�#1��fdr,op7��_����lp>oh���O�~ ߏ�d&gts���&dޏ�/`�o�o
�J?<�vrF����v.R���Ɵpld�56�%4�0/����reeK�m�XP�)�KCO*O|%56 ?�OZ� o~����E$�io����jߠ���l� ����OR��LO1Fvod��_IF��$� � ߪ�DߦX!B� U3ce��t�4 ���(M�O�5)e?Ƕ/����1?Q�D�uk �'�|����`�boto�����-���6�p�0eS ��on*��� ^�lB'����Տ_�q��_�rdk��4f�� C(ҿȿ¯ԯ�������̟�����
I���571��t�a3di39Tar��lփofk�������vP�a�@� PJ��|*��������3et�4epg���e�d�� E�5�R�I  Hw552� 747��21�pWel�R78�,� �0�ETXJ61�4��ATUP�  wmfh 5#45�p�"6�pk��VCAM  �7\awCR�I@ ED" G U�IF)!28  =j�CNREM�`��63�a�SC�H  4C D�OCV� CSU�i�!0 D s�EIOCE�54��#R694 we!!ESET=S#!3!��a 73!fanu�MASK���PRXY�_"78� �0�OCO��"�3=P[�#"�ER �J�" 7�!!J7�74#!39�  Eqq�G1�LCH 0�#OPLG%J5y000#MHCR)%sPS�17#MCS �4D"�04 O#J55< [#MDSWe!Y13MD#1s#OP#1#MPR$07�0w"0p�#�  �#PCMX �#R0A�#� &�0�0�#� ( �&0�$590( �#PRS� 3�J6903FRDz@ 02RMCNy�7ndM�93 �SNBAA�8�00�@HLB  �"Lo�SM�A0� (Ww"4 oni�t#!2  II)��TC [#TMI�Le �B�`0"K3��@TPA� �QT�Xa�t\j�@ELL�BM250`0/D8�v�$78�mon�1�95d SD95\FU�EC 0OP� UFR(@ ��;!C@ \�@;!uO�0pt"VIP�@�#� I�@0�!CS9X� �#WEB �#wHTT \stB�24 �#CG�Q#I�G�Qtopm�PP3GS!��PRC�@S#H7���w!6( �8��![�R RBB-� Ci�B01rog�w!#IF#"098`-!!` �@�A64�(AaNVD�!Ld�1h 6a68( c�`d �SR7c!te.p� 0kaч@�bc`� �CLI$0?�sb$c9�G MS�"5a�` -� A� STY�@a;l �@CTO �CwJNN0J98��ORS�0G��b�g� J�`OL�1Ab�n: SENDu�to�!L�Q���@*r#�SLM� 8�"FV�R� MCHN0CSW!SPBVP�� KPL� ds �qV$0��cCCG $p�aC�R�0
Np�QB� 8�7.f�QK� j7a0*`�p�0'3CSq7Too�CTQ��&�qTB�P�N��@In;pqC�@�Q#�� �p,#�p ��. %��$07#%� `8D#TC6� QSQ"TE� [#Xm� �tTE� gt"m�P�TTF�Q[����@�#CTG�Q�"����@�#CTH `�TT�I�@#CT'Qeqs�PCTM�@SC��$0gS��0bodyzqP�@  ���� �1� d��q�aus�a9��P�[�qW `@06; GqF `8�V@VP2@ G623R i��@j?��g� `n�g�B `"D g�D `��g�FX wmna"PVPI���+ G V�!#V	` 7 23�RVK�@Np��@CV�Q31�9�34.�vo R�erne땗��$��i��r��땁h���A���3�7� ��"�\srv����b�3b�/- Sr�B"0��<�A�J935땿B^�5 (S�O�� �g �1�1�R�|�j93땷b��E�N�5�� awm��SK� Lib �������� ����	 �"|�h��h�#��b�wmsEk�nE����q�6��pyE�  ����!�02�t Fu�ïբ6ۯm��ujKi-�I&���8k� �8!�Ń�땼P��2�2�2�Mai'�on��_�/r�;pڦh;�;�G��_r���!��4\ֶORCt��+�5�� "T¦aTP��hQ�652�a1��4���<�xk��(���ߦ�t�P��Q�rֶSB�� ch_ ����)�t!0�B�"̿ h�h땇�;���c� �����������>�<�Rp� \toֶ3�F��cl�W��2p� "���������� F����b� Qt�a�ϒ�0t��ܐFsȒ�7�6�p�t	� Ad���582��ob��|*{�\a���FMQ ���A�mcigֶ�I�or�pwI�j�rfm���Fc���@1�EYME~� w���R��b�4�K2Х70.�9E�ld,�C�6� 1PTP]��\�.�"AD.�F�p&3 k���ask�D�ȍ`4���۳dֶ�ے��ER~�7 R �ƫ/�T�?)�e�rv�G?Y?k?}?�?�?ӹapa��	d�Ъ��r�4�M��teD����79!J�d/�2��G�p�ac�T� �<6�b�/� QO��$vc>�,@Vg�����eYW��5/� 1BJ�h���R5:�d���0�@��I_��raj��e��he(}�$`��5(Xa�@���et榻�1Otdj���,�_h�\	UI�/k�jo�FO��`^�°�F��r��qW65�q���K �'6ڦus W'�b,'��'?:��n��MFR��;�]�lf�ǯ�fr>֛�w�p�/�,� �_U[ǀ�мn�x'_ i�{�����O���pJ����[@�o�in7L��O�9�\^� � R����+m�i2״h �j��҇-� f�nt >�M�A H�I  �H5529� �(Cߑ21��leR78�c�ߒ�0AcaJ6�14���0AT�UP�����545.�t-fl�6yE=��VCAM�tFLXCRId���o�wUIFULX ��28��mo�NRE�u'��63��WQ��S�CH��Cn�DOC�V�gϠCSU1�c�xr�0$�;�EIOC%tx\cF��54�oQ��9T��;�ESET�Tem!o?�S�/��7S�{�oMASK��70���PRXY�T�`��7t��`�OߐOCOe��\?�3�ô`>��0�{�?��|�-��o7n G?�39!'ߑ�õ H82L�CHd��@IOwPLG�tCGM?��0��GЎ�MHCR��Go�S�/1_�CSn4�cgm��50T�ě?�5$�[���MDSWMf.�D�����{OP��X/2L_�PR��K�����{��n�883n�CM��/0iA,��0�Ő`z~�5#�\h88� ��+�?�D���.?����4��0D�3��o�S�4����9��,i�FRDd�/2E�/��MCN5�H9y3�K�SNBA�U�"R��HLB��S�M�՛ñ�T���J512�SaߐTC4�\�TTMILe���P���A|�TPA����TPTX��5N��TEL�ԫ�0��P��8�˳���K��95����95��8�88��UECd�r;t �UFRd�_�_�Cd�2e-�VC9O4��VIP�;���I�TAX~�CSqX�����WEB4����HTT4�ka���2T�2M/So�G<#��QIG��< �.�IPGS=t\r�xO�RC��aߐ7��/a��6D�s@>�R7#��!��Oq�Ҥ� �P��Ҷ;�A���KÑ�.$�0 "��4�����NVD4���#�Ad�ap��8D���68�����R7���P��D0��a��o�bܠ. 7CLI��l\-C���CMS�'��4�wd "ްSTY�n[�CTOT�tl��sNN����ORS4ĸ;�1 ��ltiΰO	LS�( E���0�TЊ��L��6�@���9�@ ��LM4�HV� o�VR���CSshc>�PBV�4䫁/�PL�
AP�V��ust>�CC�G4��0nCR�4 H5��B���=K�H573���x?����\cms�n#�st.~TB��P�! ��7�C��x��?"�awsh?"���I0?"��3�T�Cd�K�A 4�\sl�"EĤpP��� 4�C[П"Ԥ8c��"4�(�.�CTF��c��"����CTG�73�m#G�THd�hd� �I��K�CTC�;59m�CTM�5�M����Q0��re\g�P���12�@�04�����%S��13MCTWd�9l[@_�GFd�SE]�P2d�t+��2�ա ��2d�ell��PBd�I���1Dd��a�1�F��tap VP�Id���CV�!Vtq��UA��CVK��ۣCV#�coreAL���H"�Hp!8�HK"�Hatc�J$�H�4�I� �IL0H�I�2�H��H+2�I�L�Y4=�H���Iec\a�I�2 Z93�I@{�H�@NZ+��H 1�F�K48�Z<A�Ht{@�Il �Z;"�O�Fs\! �Hk"�H{"@o�F[�PZ!o�Z���J��Tok���H��H\��Il�Z���Z2=[ng-[gToo�I�p�j(�nj�robt_�Xbt1.�JL� iur�o�I@��i�!��F��POz�ling�j��y���Y"r^zۢ�I�p��Geat^j�]��Z��_je�����_��lkҠHm,��H|��Zz��A�I  �_��  ���Gvhm��J{�svnj���H4�9\�J�@L�Ij7�49{P�Zt\j0Nj�@_"g.pjmgcal�0�fu�J��^zhm-��_bg����o�\ͫ �1�H!� j��;����MT "�(Cu�zk��&bgft�JlpX����GCT"���Gfc<]�˝26\fߟ�926�l\� Ίu��>m��;�Mul?�Q��7\^�K����7-[˝���_�61nNj48.� H- ԠH�@R_�L^ziPae��K�Я�F8\}��}�����Ћ� � R<k,�ticMoj+@�OoQxs-@�"�3�C�S j+}LB-[5s HNj+� co~��L��z��f�k˝lb�jll����-˜��k/�.���LЎ�ki;pJ/�on,�J\A���8�SK"�� ��uto�o B�������kwm� �o��Htp�ʜ n}F��ex-�˝��x��J�a^jlL�je����i��a��/����rej�1X�o�Vor�zR�ߎ��e T�Z[��[l#clN��߭�SOžgGZD��to�{�+B�H643N�`�S1G/o��sg�a�Utui��;`�J���`�;�ndm�ndiN�{/�/�/�/�/�/ �/�/??/?A?�?���riΪ! -Kj9�50/�n �zk]8c95n/�O�t �Z��wsg�K,�>��wiag� SGJ�Ю�ogu���KO�]Ltw>_@	J64t�1�s�{F O>�F�cdݛ��`3_���r-��N74�y�-�3��RINnzlly��(m^���L����sgc�zI" �#?
+�oߡ\tw /��0.�@�"���f��_�[y�Kmm�K}d�ct^�t]�+�
P�RZWCHK
kA,�;;`y<p��lK�t��LN*R85j� �@_jR ���t�iN�g WJhe�cN�L�F����wl�Z|*�dat��ʛ�greN��o�  ST�D�r7LA[NG�Aoc�e�`���Q�7��R8�70�{��8 (=P�ogge���!�58\�P�ATTs�� �t\���c "B�@Vx��1�patd���O���������{q㕔�5�a�p[�m��\㕻�7�\aw ��@�a��p6���x��ϯ�gmon���d��0�B�m�;A���\ ö��K�I�M�HCR�51 H�����g\o��@��R]� H54ۿm�<@�E���;!�����o#mm�;a��R�|�N㕬0F�C��W�P�)Ai6�� Fƫ�{�.�itx�#{ ���iaio����De�6�eve����72� R�@RƜPg��a�dl��nt��K�RBT�tOwPTN`772'�CTK"'�g�(䔠<�)� "AZ'�;q8'�q'�tzn&�{ �E'�Ama��- �Mu��ncInDPN����Ҟ��872��|�d��(��������#����masy��y �"M��o��䃲��et����\p1�����d\ ��f���lZ����lp���9���`��8+ V��ail��?� �䇢�䓢��zd�<��k`��73.f��iwrdg��- i���e\ ����� S0.j�021"�1W ��p(�`�4�� (i��e,"� "���+�^��core_�I���l`F��AY��AB���@����H�����AwBIC��Par;�M�ai������<�v c\�ITX>����  ����1���g Jcl;ib��ShiW�x4�� t994\��VSSF��� tt�\j9�f "O��w� t��$%ini�/��pٰ t�5G8�&,� t\vsR&x��L�%w� tamcl<S/+ref.�%#� tj��%m�� t[A΃&4\z�/�,z_�v�%A�%�a�%_o�l6��l% �%en	d�/<c?.?@?R5�o[?m>�6�/�dsh9f�/+trt�?<xOAE�'F  !�G0��$%��5vi�6���6 J92�F3��%O25 (�%�@e&�P�%k�4O dnw�zF��T�&`�XEpn��&g��? nw\nL�?�,nd�V��N;XfnF j���%se�V I/
&�q&фU���5r w�%/F�� �F�_�rclR&0X\pw/Y�90�Eo`t/"5Of "U//A+dprm�%g¨%��Xrsu/kmS�T_ L`�6/OŔpM�LO�j���nO1|h�ODnopn�|YCwrpR/��l���E<�Pe\ga<��Krgas�o�k���f�v��4xt�f�?m$ra�o�la`0�omk�_�TamN6�+�4�`'9K0.v �Wې�%�@�Ft��XE� sV��ДJ73=7�%|*�%,P̲�hB "+��Kwc�fF& I����99�8�vtomzFut vV�_	o;�YC��F�:8\F&�Y/� 0:��f��deb^V���$�0zFؠ"��gL���<9\�&��9�W�r}  �su"�st��G��X �f� U (�fagn�F PzFϜ6�Via�TX����vd��w��g��HzF7- O�W CH� ��$723�F���E( A�ÿտ2蚽Wc��W�svF& S�W�JRi6��_�RVo RV0���ӊ��vt�MG\etF�XoN�o�FAr��x���+�1T�F�?teR� J58��O  34	Wgl�e,�%,�j�Dq\t0"��zFwIta1lU#TA�VϜ�gw韗M�ad�W�Oa���6d� M��e�FT��9�0 H�%NT��R�69������ir�\ʆMIR��ӊenʆv���F|�3��I'TCP��Ta0�p���(MM7G�eT�o/ \tpʆI��YB'busJ׈�m��I�@zFȀ��F�����t/��W�'g, ��4`R_(!sw�&s_YC�67\JF��Tf_����Dfw��W��4gachg��a96_�d�� _���_rV��% 99�YA�e��$F�EAT_ADD �?	����~�  	�$ YA//%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /�A�S�e�w߉ߛ߭��������DEMO� N�   ��*� �2�_�V� h������������ ��%��.�[�R�d��� ��������������! *WN`��� �����& SJ\����� ���//"/O/F/ X/�/|/�/�/�/�/�/ �/???K?B?T?�? x?�?�?�?�?�?�?O OOGO>OPO}OtO�O �O�O�O�O�O___ C_:_L_y_p_�_�_�_ �_�_�_	o oo?o6o Houolo~o�o�o�o�o �o�o;2Dq hz������ �
�7�.�@�m�d�v� ������ƏЏ���� 3�*�<�i�`�r����� ��̟����/�&� 8�e�\�n��������� ȯ�����+�"�4�a� X�j���������Ŀ� ���'��0�]�T�f� �ϊϜ϶��������� #��,�Y�P�bߏ߆� �߲߼��������� (�U�L�^����� ����������$�Q� H�Z���~��������� ���� MDV �z������ 
I@Rv ������// /E/</N/{/r/�/�/ �/�/�/�/???A? 8?J?w?n?�?�?�?�? �?�?O�?O=O4OFO sOjO|O�O�O�O�O�O _�O_9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l���������Ə ����)� �2�_�V� h����������� ��%��.�[�R�d�~� ������������!� �*�W�N�`�z����� �����޿���&� S�J�\�vπϭϤ϶� ��������"�O�F� X�r�|ߩߠ߲����� �����K�B�T�n� x����������� ��G�>�P�j�t��� ���������� C:Lfp��� ���	 ?6 Hbl����� �/�/;/2/D/^/ h/�/�/�/�/�/�/? �/
?7?.?@?Z?d?�? �?�?�?�?�?�?�?O 3O*O<OVO`O�O�O�O �O�O�O�O�O_/_&_ 8_R_\_�_�_�_�_�_ �_�_�_�_+o"o4oNo Xo�o|o�o�o�o�o�o �o�o'0JT� x������� #��,�F�P�}�t��� ������������ (�B�L�y�p������� ���ܟ���$�>� H�u�l�~�������� د��� �:�D�q� h�z�������ݿԿ� �
��6�@�m�d�v� �ϚϬ��������� �2�<�i�`�rߟߖ� �����������.� 8�e�\�n������ ��������*�4�a� X�j������������� ��&0]Tf �������� ",YPb�� ������// (/U/L/^/�/�/�/�/ �/�/�/�/ ??$?Q? H?Z?�?~?�?�?�?�? �?�?�?O OMODOVO �OzO�O�O�O�O�O�O �O__I_@_R__v_��_�_�_�_�_�_m  h$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ� ����0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲�������|���  � �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p�� ����� ��$� 6�H�Z�l�~������� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ����������	�,�>�P�b� t����������� ��(�:�L�^�p��� ������������  $6HZl~�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o�i�$FEAT_�DEMOIN  �d�D`�`�,dINDEX9k�Ha�,`ILECO�MP O���zaGb'ep`�SETUP2 �Pze�b� � N �amc_AP2BCK 1Qzi?  �)h�o"�k%�o`}` Ae�om�o� � �V�z�!��E� �i�{�
���.�ÏՏ d��������*�S�� w������<�џ`��� ���+���O�a�🅯 ���8���߯n���� '�9�ȯ]�쯁���"� ��F�ۿ�|�Ϡ�5� ĿB�k�����ϳ��� T���x��߮�C��� g�y�ߝ�,���P��� �߆���?�Q���u� ���:���^���� ��)���M���Z���� ��6�����l���% 7��[��� ��D�h��i�`P��o 2�`*.cVR`� *c������JPC���� FR6:D�.�4/�TX` X/j/�U/�,;`%/�/�*.FM�/�	��/<�/<?�+STMG?q?��]?"�=+?�?�+H�?�?��7�?�?�?EO�*GIFOOyO�5eO"O4O�O�*JPG�O�O�5�O0�O�OM_�JSW_�_�� Sn_+_%
J�avaScript�_�OCS�_o�6��_�_ %Cas�cading S�tyle She�ets0o� 
AR�GNAME.DT_o��0\so1o�Q�d�o`o�`DISP*�o�o�0�o7�e�)q8�o
TPEI?NS.XMLg�:\{9�aCus�tom Tool�bar��iPAS�SWORD.��FRS:\�� �%Passwo�rd Config@���������� �r�����=�̏a� s����&���J�\�� ������K�ڟo��� ����4�ɯX������ #���G�֯�}���� 0���׿f������1� ��U��yϋ�ϯ�>� ��b�t�	ߘ�-߼�&� c��χ�߽߫�L��� p����;���_���  ��$��H����~� ���7�I���m���� ��2���V���z���! ��E��>{
�. ��d��/� S�w�<� `�/�+/�O/a/ ��//�/�/J/�/n/ ?�/�/9?�/]?�/V? �?"?�?F?�?�?|?O �?5OGO�?kO�?�OO 0O�OTO�OxO�O_�O C_�Og_y__�_,_�_ �_b_�_�_o�_�_Qo �_uoono�o:o�o^o �o�o)�oM_�o ��6H�l� ��7��[�����  ���D�ُ�z���� 3�ԏi�������� ßR��v�����A� Пe�w����*���N��`���֦�$FIL�E_DGBCK �1Q������ ( ��)
SUMMA�RY.DG�����MD:3�s����Diag Sum�maryt���
C?ONSLOGi�L��^�������Con�sole log�����	TPACC�N�R�%:�wς��TP Accou�ntinρ�F�R6:IPKDM�P.ZIP�ϯ�
����σ���Exception ߱�_��MEMCHECK�m�Կb����Me�mory Dat�a��֦LN�)n�RIPE�\�n����%�� Packet L�κ��$SA���ST�AT�����ߋ� �%�Stat�us��<�	FTP�����r�����m�ment TBD���� =�)E?THERNEU����B�S�����Eth�ern(��fig�ura߇���DCSVRF���������� veri?fy all٣�M(��DIF�F����/d�iff�PB���CHGD1�x�� �FQ&���	2�� q5�YGD3�8��'/ �N/��UPDATE�S.m S/��FR�S:\k/�-��U�pdates L�ist�/��PSRBWLD.CM�/«��"�/�/�PS�_ROBOWEL<1���:GIG�ߊ?�/�?��GigE� ��nostic�*�ܢN�>�)>�1HADOW�?�?��?5O��Shad�ow Changye��٤&8+�2NOTI��O"O�O���Notifi�c��\O٥O�A ��_��2_կ?_h_�� �__�_�_Q_�_u_
o o�_@o�_dovoo�o )o�oMo�o�o�o�o <N�or��7 �[���&��J� �W������3�ȏڏ i�����"�4�ÏX�� |������A�֟e�� ���0���T�f����� �����O��s��� ��>�ͯb��o���'� ��K��򿁿ϥ�:� L�ۿp����Ϧ�5��� Y���}���$߳�H��� l�~�ߢ�1�����g� �ߋ� �2���V���z� 	���?���c���
� ��.���R�d�����������$FILE�_� PR� �����������MDONLY� 1Q���� �
 �)�@_V�DAEXTP.Z�ZZ��p�G�L6�%NO Back file !��U3�M��7 ����G�&�J \����E� i�/�4/�X/� e/�//�/A/�/�/w/ ?�/0?B?�/f?�/�? �?+?�?O?�?s?�?O �?>O�?bOtOO�O'O �O�O]O�O�O_(_��?VISBCK����>*.VD)_s_��@FR:\BPI�ON\DATA\�^_R�@Vis?ion VDt�_ �O�_�__o_Ao�_ Rowoo�o*o�o�o`o �o�o�o�oO�os �@�8�\�� �'��K�]����� ��4�F�ۏj����̏ 5�ďY��j������ B�ן�x����1����ҟg���MR2_G�RP 1R���C4  B�O��	 
������E��� ֯�r���O�HcEP]��O��#M��
�/KA���?�&��r���:6:N{�R�9-�Z���A�  v���B�H��C`}dC�{�N��B�{���r���пὫ�@UUT��U����/����>��>c���>rа=ȫ��>i�=����>����:���:��:�/:6)�:��~ϗ�2ϔ��ϸ�������z�_CFG {S��T  ��a�s߅�0[NO ���
F0�� ���/\RM_CHK�TYP  ����O����������OM���_MIN��L�������X��S�SB7�T�� ��5�L�,�U�g����TP_DEF_�OW��L�����I�RCOM�Ѝ��$�GENOVRD_�DO��	��TH�R�� d��d��_�ENB�� ��R�AVC��U�UQ �Υm�X��|��q������ � �kOU��[��O�����⾥8��:���
,.  C�x �h�������B�ϡ�����\n�!�SMT'�\.����+�w�$HOS�TC7�1]K[s�Y��� MCL���MI� _ 27.0�1�  e}���  /*�1/C/U/g/��!/#	anonymous�/�/�/�/D�/? L��8; {}/j?��?�?�?�? �?/�?OO0OS?�? �/xO�O�O�O�O?UO +?=?_QOs?1_b_t_ �_�_�?�_�_�_�_o '_]OoOLo^opo�o�o �O�O�O_o G_$ 6HZl�_��� ���o1o� �2�D� V�h��o�o�o���ԏ ��
��.�uR�d� v�������?����� ��*�q��������� ��ݏ��̯ޯ��I� &�8�J�\�n���ǟٟ ��ȿڿ���E�W�i� F�}�jϱ��Ϡϲ��� ��������0�S�T� ��xߊߜ߮����� +�=�?��s�P�b�t� ����ϼ�������� '�]�o�L�^�p������/ENT 1^��� P!���  ������* ��Nr5~Y� �����8� \1�U�y� ����4/�X// |/?/�/c/�/�/�/�/ �/?�/B??N?)?w? �?_?�?�?�?�?O�? ,O�?ObO%O�OIO�O�mJQUICC0 �O�O�O_�D1_�O�OV_�D2W_3_E_�_�!ROUTER�_�_�_�_!PC�JOG�_�_!�192.168.�0.10�O�CCA�MPRTGo#o!b7e1@`noUfRT�_�ro�o�o��NAME� !��!RO�BO`o�oS_CF�G 1]�� ��Auto�-started^��FTP��~q ���F����� ���9�K�]�o���� &���ɏۏ�����W i{X����o����� ğ֟������0�B� e��x���������ү �������Q�>���b� t�������q�ο�� ��9���L�^�pς� �Ϧ�������%�� Y�6�H�Z�l�3ϐߢ� ��������}��� �2� D�V�h���������� �����
��.�@�� d�v���������Q��� ��*<���� ��������� ���8J\n�� %�����EW i{}O/��/�/�/ �/�/��/??0?B? e/�/x?�?�?�?�?�? /+/=/�?Q?>O�/bO tO�O�O�Oq?�O�O�O _'O(_�OL_^_p_�_��_(�`_ERR �_z�_�VPDU�SIZ  9P^�S@��T>�UWR�D ?EuA� � guest3V$o6oHoZolo�~o�dSCD_GR�OUP 3`E| uIq?YM �nwCON�nTAS�n�L��nAXP�n_E��o9P�n�RTTP�_AUTH 1a��[ <!iPendan�g�~@}�9PJ�!KAR�EL:*���}�KC����pV�ISION SE!T�`E��I�!\�J� t��s����������Ώ���-���dtCTR/L b�]~�9Q�
`�FFF�9E39�DFR�S:DEFAUL�T��FANU�C Web Server����bvo dL��'�9�K�]�o��TWR_�`FIGw c�e�R����QIDL_C_PU_PC9QsB�@� BHǥ�MINҬ�a�GNR_IO�Q�R9P�X�ɠNPT_SIM�_DO�!�STAL_SCRN�� �y�+�TPMODNTOLY�!���RTY8��&�9�hp�ENBY��cƣO�LNK 1d�[ �`�����1�C�UϾͲMASTE����&�OSLAVE� e�_˴jqO_gCFGsϦ�UOD�|�Ϩ�CYCLE����ļ�_ASG 19f���Q
 W�9� K�]�o߁ߓߥ߷��߀�������#�_��N�UM�S�b�U
��I�PCH��j�O_R?TRY_CN�x�Z��U�_UPD�S����U �������g�θ`��`ɠP_�MEMBERS �2h��` $�e��>��HyɠSD�T_ISOLC � ���r�\J2/3_DS��q���?OBPROC��%��JOG�d1i���89Pd8�#?�.���.�?�?�?OQNs��V����3W~�����������POSR�E��$�KANJI�_m�K�i�pMO�N j�k~�9Ry ����//�^�r��k����9%Th���p_L�I�l�kEYLOGGIN����`����U�$�LANGUAGE� ����� ,�!�QLG��lq�9R마9Px�p�  ���砬9P'0�3X�k���MC�:\RSCH\0�0\��� N_DISP m��DA8MK�SLOCw�آ�Dz ��A�#OGBOOK nۄ��9P~��1�1�0X�9O%O7OIO[OmN`�Mɱ���I��	�5@Ib�5�O�O�5�2�_BUFF 1oؽ�O2A5!_�2 ��=_?7Y_k_�_�_�_ �_�_�_o�_o:o1o CoUogo�o�o�o�oe4~��DCS q�= =��͏L�O-��1CUg���bIOw 1r� ���s20����� ���1�A�S�e�y� ��������я���	���+�=�Q�|uE�TMl�d����Ο�� ���(�:�L�^�p� ��������ʯܯ� �8��7�SEV��u=]{�TYPl���`z�����!�PRS����/S��FL 1s�}����$�6�`H�Z�l�~ϯ�TP� �l�i��=NGNA�M��A5�"e4UPSFm0GI��\!�����_LOAD��G �%u:%CON�ROD4U9�:�MA?XUALRMI�c�8W�T���_PR�����3�R�Cp0t��9�M���3Eݗ���Pw 2u�� �1V�	i�00��� �߭�1��.�g�x U���������� ���8�J�-�n�Y��� u�����������" F1jM_�� �����	B %7xc���� ���/�/P/;/ t/_/�/�/�/�/�/�/ �/�/(??L?7?p?�? e?�?�?�?�?�? O�? $OOHOZO=O~OiO�O�K�D_LDXDI�SA����zsMEM�O_AP��E ?=��
 b��I �O_"_4_F_X_j_|_~R�ISC 1v�� ��O�_ ���_��_�Ooo@o�_C_MSTR w:�~_eSCD 1x�M�4o�o0o�o�o�o�o P;t_� �������� :�%�^�I���m���� ��܏Ǐ ��$��4� Z�E�~�i�����Ɵ�� �՟� ��D�/�h� S���w���¯���ѯ 
���.��R�=�O��� s�����п����߿� *��N�9�r�]ϖρ����PoMKCFG �ynm����LTAWRM_��z����и���6�>�s�M�ETPU�ӫІ��viND��ADCO�LXի�c�CMNT�y� l�g` {�nn��-�&�����l�P�OSCF����PgRPM����STw�{1|�[ 4@�P<#�
g��g�w� ��c��������� ����G�)�;�}�_��q�����������l�S�ING_CHK � |�$MODA�Q�}�σW��#D�EV 	�Z	�MC:WHSIZ�E�M�P�#TAS�K %�Z%$1�23456789� ��!TRIGW 1~�]l�U%�\�!�S
K.�S�Y�P�69"EM_INF 1�� `)�AT&FV0E�0X�)�E0�V1&A3&B1�&D2&S0&C�1S0=�)A#TZ�#/
$H'/O/�Cw/(A/�/b/�/�/�/? �&?� ��/�?3/�?�/�? �?�/�?�?"O4OOXO ??�OA?S?e?�O�? �?_CO0_�O�?f_!_ �_q_�_�_sO�_�O�O �O�O>o�Obo�_so�o K_�owo�o�o�o�_ �_L�_o#o��Yo ����o$��H� /�l�~�1��Ugy ���� �2�i�V�	��z�5�������ԟPN�ITOR��G ?�k   	EOXEC1���2�3�4�5�� �U7�8�9��� �������(���4��� @���L���X���d���Pp���|���2��2��U2��2��2��2ŨU2Ѩ2ݨ2�2���3��3��3(�#R�_GRP_SV �1�� (�ſ1x�>Ka����|�ӣRƮ_Ds����PL�_NAME !����!De�fault Pe�rsonalit�y (from �FD) ��RR2��� 1�L6(�L?����	l d��nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲�����B2]���*�<�N�@`�r����<�� ��������,�>�P��b�t�����BJ�  �\  ��  ������  A�  B���T��� 
��������  �������B��p��ȷ  CH CH P� Ez  E��� E�` E��;%�Z��*� �  Ec��F�@&���T Ai�  dx�H�x�	@$Hxd�dڭ�}`(d�� 8(xx$$Ay Xtd D (DDdpWwX ��	X�vXHXH���/y�y 	(� !��  7%3E	��Em�X�w$%XH$%P�� �/�/�/�/�/�/?�?+?=?O?a?s=F��r?�?�?�?�6���E�2ExB�2�������?K
زd��'O9NO\O�jG�0��|M��ն'�4 � Wq%�O�O�N �0h�G�O�JA  A��C����_�OC_9W�  � TB�LY��
��_�\��Q�Y=²CÈ�V�`HR0� ʒ�P( @7%?���a�Q?ذaر@��6�&س��2n;��	lb	 � ����pX��U�M`��X � � ��, �rb��K��l,K���K���2KI+�KG0�K �U�L�2o�E	O�n��@�6@ t�@?�X@I��b`��o�C�N�����
��}v��G���` q�m�|�~kQ�
=ô���  Hq�o`!b��s�  ���a�  �����ذa�s�G��d�}�m��o�q��v��O��E	'� �� 0�I� ��  � Q�J:��ÈT�È=�s��l���@|�@��}~�Q����R��Ȼ��N8���  �'��ap?�ɡ�b!p�b){�B��?�CIpB  X��=ذ��C�A�g!	���o�P�IB P���8�����P��ԕرD  �O���O��A�,�:��Š
�`l�1�	 ٠p�*�� p` l`:�4�  �t�?�faf{O��įV� �P������a�!�/�?Y�)R�a4�(ذ]�P�f����a\c\dƃ?3�33-d���;�x�5;��0;�i�;�du;�t�<!�+}�oݯ���b�Sb�P?ff�f?��?&�9�@��A#$�@�o[,ž�x�	� &f6�ed�g���Hd 㯸ϣ����� ���$߀�H�Z�E�~߾�&eF��mߺ�i���U��߰y���2���E�0 ����y�d������ ��������?�*�܏ r�8�.o�ߺ����T� );ڿPb�� ������P��cA��T C�`=�ϵ��Y}��2��������C���W�C�= �` #Ca��������(!�`�<���bC�@_;C9�B�A�Q�>�V{È�����Y�uü��
/���Q���hQ�A��B=�
?h��Ä/iP��W���ÈK�B/�
=�������=�K�=�J�6XK�r#H��Y
H}��A��1�L�j�LK����H:��HK���/0	bL ��2J��8H���H+UZBu�a?�/^?�?�?�? �?�?�?O�?O9O$O ]OHO�OlO�O�O�O�O �O�O�O#__G_2_k_ V_{_�_�_�_�_�_�_ o�_1oo.ogoRo�o vo�o�o�o�o�o	�o -Q<u`�� �������;��&�K�q�\�����G�y����� C�a>ɏ Ĉ����OCVF�����+<b����Kc�f�� 
E����T�ٟz�(��_�h۟攱�����N��������3lC�8(�:�H���T�f���t�.3��}�����k���q'�3�JJ�����@گ���4�"�]P̲	Pf�������⟛�0ſ���Ի�����/��?�{?�N�u�  fUh�*ϳϞ��� ���Ϣ�t�.��R�@ۃ�X�bߘ߆ߨ�)�Z�ߺ�  ( 5�	������B��0�f�t�  2 wE%p"E[@��N�"BC%��%@ߏ�� %������)�;�������������%(n�n�%��%r��Xc
 �� !3EWi{�� �����b*[���P�I�v��$MSKCFMA�P  ��� ^�����p�DONREL  �X�[��DE�XCFENB�
8Y�FNC���JOGOVLIMҍd��dDKE�Y��%_P�AN�""DRU�N��>#SFSPDTYw�����SIGN��T1�MOT��D_�CE_GRP 1-���[\���/ ��?&?��?Q??u? ,?j?�?b?�?�?�?O �?)O;O�?_OO�O�O LO�OpO�O�O�O_%_ _I_ _m__f_�_O��DQZ_EDIT��$UTCOM_�CFG 1�Q��_o"o
�Q_A�RC_�X��T_MN_MOD����$�UAP_�CPLFo�NOCHECK ?Q W����o�o �o�o'9K]�o�����vN�O_WAIT_L؉'�W� NT�Q��Q���_ERR��!2�Q���  �_t�������*���Ώ�d``OI��P�x� 3搓_���8�?��4����|�B�PARAMJ��Q���	������s�� =��345678901�� � ���?�Q�-�]������u���ϯ����������7�ODR�DSPEc�&�OF�FSET_CAR8�PKom�DISz�K��PEN_FILE����!$a�V<`OPT?ION_IO
/=!�аM_PRG %Q%$*	�ά�WORK ��'=� ��K�7:U�h� ���f�9(�f�	 ���f��5���M�RG_DSBL  Q�����L�RIE�NTTO* ��C���Z��M�UT__SIM_DطX�+M�VQ�LCT �%��R_�$aQ�'ԏ_PEXh`��b�R[AThg d�b�>r�UP �5� � ����߼������$��2�#�L�6(L?��	l d'�O�a�s� ������������ �'�9�K�]�o���������H�2>����� /ASew�N�<��������1CUgyH����P�� �  ��  �U�?A�  B��P[B����H���  ���U�B��p�������N�P Ez  �E�� E�` �E��;(�����Z�/��� � E��''����@#���T�AJ(��E!Y!a!)!m! Y!u)%)!Y!E!�%E!ڎ$�^$A!�	!E! a!�%%	-Y!Y%�-58�Z 99U%E!�	D!	$D%%E!Q481 X291�%�)95�/W#95 )%91m5a!�5/Z7�%�Z (�8�1�<a1� EE	�(�Em �494X6E9=)%E15�� |O�O�O�O�O �O�O�O__0_B_T]F�S_y_�_�_�Vh�����_�[��%�on�_=oKg�]�]�&�'4 �� W%po�oX� ����g�o�jA�A=��c�����o�oT$w���tB�@(~�`��r�|�� q�y�$�O��1�'k�'��3�{`��0���P( @PED�D��q?Q�Cl��pF~��o  ;�	�lD�	u� ����pX��[�2��X � � �,i��X��`H��9H��H��H`��H^yH�R�l���_�����`�C#�B� C48ӄlŎ��9��_�
=���� �������cBz���Βa�m�另b�s�� �q����g䟒�챏Ǒ��ٖ�o���e	'�� � �I� �  �q<�=���9�K���@a�g�b����������唠����N��  '۰��Ɓ"�B�Ղ��т6���� �  ��	C�a��	m�~��p=�Bp��Н����px����D��o޿�oϰ�&��o�5�Ю�`Q��	 S٠U�f� U� Q��:���#����?��ff\o�ϩ�;� !�p����"�8� ߖ�?Y
r��q=�(� B�PK�fɆ�A�A�^��?333��m��;�x5;��0�;�i;�du�;�t�<!��y������t���r�p�?fff?x�?&����@��A{#	�@�o[� �	]������uI��w h���-��ϝ����� ����	���-�?�*�c� u�L�������4�V�X�X����EjPf� ��^I�m�� �� �$��W �������9� �/ /��5/G/�z/�e/�/�/�/�/�`�A1��$�t�/ C�/"?p�(d��>�?��P�n?�/�?}?��(���W�?C�@�` !CT��?�j4�j0i1�A@I�!����bC@_;C9��BA�Q��>V`.È�����Y�u�ü��
�?�3���Q��hQ�A��B=�
?�h��iOJp���W��ÈK��B/
=�����Ɗ=�=K�=��J6XK�r�#H�Y
H}���A�1�=L��jLK����H:��HK��O�@	bL� �2J��8H���H+UZBu�?F_�OC_|_ g_�_�_�_�_�_�_�_ o	oBo-ofoQo�ouo �o�o�o�o�o�o, P;`�q�� �������L� 7�p�[��������ȏ �ُ���6�!�Z�E� ~�i�{�����؟ß�� � ��0�V�A�z�e��Gϭ���� C��a�/�� Ĉ��<ЯׯCVF������üKG�j���K<H�K�� 
Ep�s��9���90(91�_ʙh��y����i���N����T�3l�C���-¢��9�Kϰt�.3��}e�w�k���q'�3�JJ�� ���Ͽ�������B5%P��PK�Zgt��ǿ�ߪߕ��߹�� �������$�{$�3�Z�  fUM��� �������Y��7�%��=�G�}�k���)Z����  ( 5�� �������'KY  2� E%pIFE[-@tN�IFB�!�!�� C��0� T�@ į����*H3��Tfx��PT�T�94���T�D=4H;
  �//*/</N/`/r/ �/�/�/�/�/�/�/GJ�@2��5�I�v��$PARAM_MENU ?����  �DEFPU�LS��	WAI�TTMOUTT;�RCVg? S�HELL_WRK�.$CUR_ST�YL���<OP9T��?PTB�?�2�C�?R_DECSN_0<�L	OO-OVO QOcOuO�O�O�O�O�O��O�O_._)1SSR�EL_ID  ��Y�=UUSE_PROG %8:q%*_�_>SCCRk0�ORY@3�W_HOSoT !8:!�T�_�ZT\Ю_ c�_�Q�c<o�[_TIM�Ei2OV�U)0GD�EBUGMP8;>SG�INP_FLMS�`�gn�hTR�o�gP+GA�` �lC�k�CH�o�hTYPE
5<A)_#_Y� }������� ��1�Z�U�g�y��� ����������	�2� -�?�Q�z�u�����ཟϟ�
��eWOR�D ?	8;
 �	PR�`U�MsAI@��SU�1�E�TE#`U��	�4R�COLS�n����vTRACECToL 1���B1w I�7 8��W d�ެ��DT �Q����РD� � *�Q����W .��.��.��`.��U"��	�
�U��2�:��B�B���"�2��;��3�:�B�J��+� =�O�a�s��������� Ϳ߾��K�a��[Ñ� �ϲ�����9����� ��	��-�?�̨ߺ� ����P�b�L�~ߐؓ� ��)�;��'�Y�k� }�oρϛ������� ����+�=�O�a�s� �������������� '9K]o�0 \n������ ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �uX����� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ� ���ߚ������0� B�T�f�x������ ��������,�>�P� b�t������������� ��(:L^p �������  $6HZl~� ������/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?�?�?�?�?��?�?OA�$PG�TRACELEN�  A  �_�@�$F�_UP �����SA[@?A�T@$A_CFG M�SE=CAT@��D�D�O�G6@�O�hBDEFSPD ��sLA6@��$@H_CONFI�G �SE;C U@@dT�3B AQP�D�A1Q�@�$@INk@T�RL �sM�A8l�EFQPE�E�W��SA�DQ�IL�IDlC�sM	�TG_RP 1�Yb@�lAC%  ���l�AA��;H��N��R���A�!PD	� a3C	�\T�Ai)iQP� 	 �O4VGg�Co ´|c^oGkB `�a�opo�o�o�o�o��b"�Bz��o7I~3 <}��<�oN�J �����f�)� �9�_�J�`z����@
t���d�ŏ�֏ ���3��W�B�{�f��x�����՟�����J)�@)
V7.1�0beta1�F� @�@�?�A&ff�Q2��CPC�`�D�D�k`[�C�T��@� DĠ Dr�- �QBH�`�L��P�C5R A?� � ��CCx����b���P!P��A����Ap�B�b!PA1�������
�?L��?333A@��"���Fff.��b�w.:�7��AeC�Q�KNOW_M  ��E{F�TSV �Z(R�C���� ��ʿ��ٿ�$�A�!m�SM�S�[ ��B�	�E��C�Ϗ�̓E`��2�E@�2������Z�� L�MR�S�Y�%T�j���AC5�����e@�Rۚ]ST�Q1� 1�SK
 4�U��A�¨߰E��*� �߽�������J�)� ;�M�_�q����� �������F�%�7�|���Ep�2{���A�#<�����P3��������p�4��+�p�5HZl~p�6 ����p�7� $p�8ASewnp�MAD0F [F�p�OVLD  �SK�ϼOr�PAR?NUM  /�O�//T_SCH� �[E
}'F!�)=C�%U�PDF/X)�/3Tp�_CMP_O�0@T@@�'{E�$ER_CHK5yH!6
?;�RS�]��Q_MO��o?�5_k?��_R/ES_GzФ~ݍ� �?�OO�?%OO*O[O NOOrO�O�O�O�O�O �O��3���<�?_ �5��(_G_L_�3G g_ �_�_�3� �_�_�_�3 � �_o	o�3@$oCo�Ho�3�co�o�o�2V� 1�~կ1e�@�c?��2THR_�INR�0�!7³5d��fMASS Z�wMN5sMON�_QUEUE a�~�f��0�� �4N0UH1NEv6;�p�END�q�?�yEX1E��u� BE�p�>�sOPTIO�w�;��pPROGRAM7 %hz%�p�o�l/�rTASK_I���~OCFG �h/\���DATuARè��@��2�����#�5�G�� k�}�������^�ן�x�����INFOR��܍�wtȟe�w��� ������ѯ����� +�=�O�a�s�������л�Ϳ(�4��܌ ��I��� K_���8��T��ENB� ͠�1>ƽ�I��G��2��� P(O8�ҡϳ� ������_EDIT ᭘��ߋ�WER�FL�x�cm�RGA�DJ �8�A���i�?�0t�
qLֈq����5�s?�!��<@��*�%���@�#ߊ�챳2���F�	Hpl��G�b��>���A�d�t$I��*X�/Z� **: c�0V�h���Ǟ���B����������� ���������b��� L�B�T���x������� ��:����$,� Pb����� ��~(:h^ p������V/  //@/6/H/�/l/~/ �/�/�/.?�/�/??  ?�?D?V?�?z?�?O �?�?�?�?�?rOO.O \OROdO�O�O�O�O�O �OJ_�O_4_*_<_�_ `_r_�_�_�_"o�_�_ooo�f	���o�p �o�o�dJ��oL��o#�oGY��PREF� ����p�p
~L�IORITY�����P�MPDSP�>ߴwUTz�4�K��ODUCTw��8�\�OG�_�TG;�|����rTO�ENT 1���� (!AF_I�NE�pp�{�!�tcp{���!�ud��ˎ!iccm�����rXY�������q)� 0p�/�A��p�)�j� M�Y���}�������� ן���8�J�1�n�U�$����*�s�Ӷ}}��x���,�>�%�jf�p�/z�֯K�,�������A��,  �p�������ʿ�u"�ut�}�sF�P��PORT_NUM��s�p�P�_CARTREP�p|��|�SKSTA�w� K�LGSm�͸������pUnothingϿ������c{t�TEM�P ����ke���_a_seiban0C�,S�y�d� �߈��߬�����	��� �?�*�c�N��r�� ����������)�� M�8�q�\�n������� ��������#I4 mX�|�������3��VER�SI�p �d �disable�d>SAVE ���	2600/H721:&��!;���̏� 	�(�rmoN+E/`�e@b/�/�/�/�/�*z,D�? %`���_-�W 1���E0��b8eO?a?4gnpUR?GE_ENB3��vl�u�WF�0DO�v���vWi��4�q*�W�RUP_DELA�Y �CΡ5R_?HOT %�f�q�:�.O�5R_NORMALH
�OrOAGSEMIQOwO�Olq_QSKIP-3���>3x$�O _1_C_ ]&ot_b_�_�_�_�_ �_�_�_o(o:o o^o Lo�o�o�olo�o�o�o  $�oH6X~ ��h����� ��D�2�h�z�����$RBTIF�4�G�RCVTMOU�\�����DC�R-3��I ��QE=U4�1D�͛�C�JA?͜6�ט]����q�6���1B�AY����_V�R_� ;�x5;���0;�i;��du;�t�<!���h��R���̝ �����&�8�J�\��n����������RD�IO_TYPE � 4=��¯EFP�OS1 1�C�
 x/:�H2��b�M� ��/��E�οi�˿� ��(�ÿL��pς�� /�i��ϵ��ω�߭� 6���3�l�ߐ�+ߴ� O����߅ߗ���2�� V���z���9���� o�������@�R������9��������OS/2 1��;+�u����-��Q���3 1�����G��|�gS4 1�~����ZE~�S5 1�%7q���/�S6 1Ũ��/�/o/�/>&/S7 1�=/O/�a/�/??=?�/S8 1��/�/�/0?�?��?�?P?SMASK 1�߯ )�OFN�7XNOܯFUO<_C�MOTE����X4uA_CFG ��|M�1\A�PL_�RANGxA���AO�WER ����@�FSM_DRY�PRG %�%�y?!_�ETART ���N/ZUME_�PRO�O_�_X4_�EXEC_ENB�  ����GSP�DdP�P�X���VTD�B�_�ZRM�_�XI�A_OPTION�φ����pAINGoVERS.a��z_�)I_AIoRPUR�@ @O\�o�=MT_�0T�@�zO��OBOT__ISOLC=N�F��1�a�eNAME�Rl�bo�:OB_O�RD_NUM ?��H�aH�721  V1;wLqr�qrV0.qr��sps�u�\@��PC_TIM�Ė��x��S23�2�B1����aL�TEACH PENDAN΀�7\H���x?c�Ma�intenanc�e ConsV2��#�"�_�No Use��N��r����������С�rNPQO>P�r\A<e�qoCH_LgP�|N�w�	<��!U�D1:b�	�R�0VgAILRq2e��u�pASR  ��:a�B�R_INoTVAL1f��I��+n��V_DAT�A_GRP 2�X��qs0DҐP�? `��?��o�������� կï�����-�/� A�w�e���������� ѿ���=�+�a�O� ��sϕϗϩ������ ��'��K�9�[߁�o� �ߓ��߷��������� �G�5�k�Y��}�� �����������1�� U�C�e�g�y������� ������	+Q?�uDA�$SAF_DO_PULS�p�E@�C�� CANd�r1f�vpSC�@��'�'�}��QV0D�D�qL�L�+AV2 y�'9K] o��������ڈ��2$($Md($C!u�1#
) @�Co/�/�/ȥ.W)k/ M��$_�_ @݃T:`��/??&?39T D��3?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O֏��i%�O�O�O܉x�!L� �;�o݄��p�M
�t��Dipp�L��J?� � ��jL� ��j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt ���������(�:����/c�u� ��������Ϗ��B� %�1�C�U�g�y���@������Ƒ��0R MS�EW]�$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ�����M���*� <�N�`�r߄ߖߨ�� ��������&�8�J� \�ǟ���������� ��������,�>�P� b�p������������� ��%7I[m ��������!3EWit�OB3t���� �////A/S/e/w/@�/�/�/�/�/�*���/?6��\R�?�M	1234�5678XRh!?B!̺����?�?�?�? �?�?�?OOA�>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ o]-O�_�_�_�_�_�_ �_o"o4oFoXojo|op�o�o�oq_BH�o �o�o!3EWi {�������<�v[;�j�A� S�e�w���������я �����+�=�O�a�xYD�k�������ɟ ۟����#�5�G�Y� k�}�������v_ׯ� ����1�C�U�g�y� ��������ӿ���	� ȯ-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�σߕߧ߹� ��������%�7�I�[�m�����v6����z��!�3��O:Cz  Aоz   �@�2��v0� @�
~���  	�r�������������ph�u�����K] o������� �#5GYk} ��0����/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-?�G�������*@  <�X4t��$SCR_�GRP 1�'�� '�� t� �t� �E5	 �1��2�2�4�� W1G3�;97�7�?�?O�C��|�BD�` D��3NGK�)R-200�0iC/165F 567890���E��RC65� �@�
123I4�E�6t�A�����C�1F�1�3�1�)�1A�:�1�I	���?_Q_c_u_�_���H��0 T�7�2�_�?�_�_o�6�t��_Lo�_poB8�boK�h�@�UO���eBǙ�B��  B�33B� �`�e�b�c�1Ag��oG  @t��e�1@>@�	  ?�w�bH�`2�j�1F@ F�`\rd[o�s �������*� �9�a�a)rU�@�R�d�v�B����ʏ��� ُ����H�3�l�W� ��{���Ě2C�?���7���9�t�!q@"p>SԪD_�U��r�`y��`ȏ�@�G�L�3��ϯ�A>G��1��"oe��)�t� �<�N�\�*��q�}���^� P���(����ӿ�g1E�L_DEFAUL�T  �D���t���HO�TSTR� ��M�IPOWERFL�  K����?�W�FDO� S�R�VENT 1�����P0� L!�DUM_EIP�翬��j!AF�_INE��ϵ!'FT�������9!�_B� ��i��!RPC_MAINj�LغXߵ�|�'VIS��Kٻ���o!TP��PU����d��M�!
PM�ON_PROXYN��e<���g���f����!RDMO_SRV���g��1�!R�DM���h, �}�!
~�M����il���!RLScYN�@����8��>!ROS��<��4a!
CE>�MTCOMb���kP�!	vCO�NS���l��!}vWASRC ����m�E!vUSBF��n4�0� �����/�'/��K//o/�RVI�CE_KL ?%��� (%SVCPRG1v/�*�%2�/�/� 3�/�/� 4??� 56?;?� 6^?c?� 7�?�?� H\��?L19�?�;�$ H�O�!�/+O�!�/SO �! ?{O�!(?�O�!P? �O�!x?�O�!�?_�! �?C_�!�?k_�!O�_ �!AO�_�!iO�_�!�O o�!�O3o�!�O[o�! 	_�o�!1_�o�!Y_�o �!�_�o�!�_{/�"�  �/� F�E1��� �����
�C�U� @�y�d���������� Џ����?�*�c�N� ��r��������̟� �)��M�8�_���n� ����˯���گ�%� �I�4�m�X���|������ǿ�ֿρ*_D�EV ���oMC:�H'�?GRP 2ׇ�+p�� bx 	�/ 
 ,y�ϒ� +r~ϻϢ�������� ��9� �]�o�Vߓ�z� ���߰������#�z� G���k�}�d����� ����������U� <�y�`���������*� ��	��-QcJ �n����� �;"_FX� �������/� /I/0/m/T/�/�/�/ �/�/�/�/�/!??E? W?�{?2?�?�?�?�? �?�?O�?/OOSO:O LO�OpO�O�O�O�O�O _^?�O=_�Oa_H_�_ �_~_�_�_�_�_�_o �_9oKo2oooVo�ozo �o�o _�o�o�o#
 G.@}d��� �����1��U� <�y����o��f�ӏ� ̏	���-�?�&�c�J� ��n��������ȟ� ���;���0�q�(��� |���˯���֯�%� �I�0�m��f������ǿ������R�d ��	�4��X�C�|�gϠϯ�%�����R������������ ���+��O�=�s߁� �Ϧ���i��������� �	��Q��x��A� �����������Y� �P���)���q����� ������1�U���I ��Ym���	 �-�!E3U {i����� �//A///Q/w/� �/�g/�/�/�/�/? ?=?/d?v?-?O?)? �?�?�?�?�?OW?<O {?OoO]OO�O�O�O �O�O/O_SO�OG_5_ k_Y_{_}_�_�__�_ +_�_ooCo1ogoUo wo�_�_�oo�o�o�o 	?-c�o��o S�O����� ;�}b��+������� ��ɏ�ݏ�U�:�y� �m�[��������ş �-��Q�۟E�3�i� W���{����دꯡ� ï���A�/�e�S��� ˯���y��ѿ��� �=�+�aϣ���ǿQ� �ϩ����������9� {�`ߟ�)ߓ߁߷ߥ� ������A�g�8�w�� k�Y��}������ ��=���1���A�g�U� ��y����������	 ��-=cQ��� ���w���) 9_���O� ���/�%/gL/ ^//7///�/�/�/ �/�/?/$?c/�/W?E? g?i?{?�?�?�??�? ;?�?/OOSOAOcOeO wO�O�?�OO�O_�O +__O_=___�O�O�_ �O�_�_�_o�_'oo Ko�_ro�_;o�o7o�o �o�o�o�o#eoJ�o }k����� �="�a�U�C�y� g�������ӏ���9� Ï-��Q�?�u�c��� ۏ��ҟ�������)� �M�;�q�����ןa� ˯��ۯݯ�%��I� ��p���9�����ǿ�� ׿ٿ�!�c�Hχ�� {�iϟύ��ϱ���)� O� �_���S�A�w�e� �߉߿����%߯�� ��)�O�=�s�a���� ���߇�������%� K�9�o������_��� ��������!G�� n��7����� �O4F�� g�����'/ K�?/-/O/Q/c/�/ �/�/��/#/�/?? ;?)?K?M?_?�?�/�? �/�?�?�?OO7O%O GO�?�?�O�?mO�O�O �O�O_�O3_uOZ_�O #_�__�_�_�_�_�_ oM_2oq_�_eoSo�o wo�o�o�o�o%o
Io �o=+aO�s� ��o�!���9� '�]�K��������q� ��m�ۏ���5�#�Y� ������I�����ßş ן���1�s�X���!� ��y���������ӯ	� K�0�o���c�Q���u� �������7��G�� ;�)�_�Mσ�qϧ�� ��ϗ�ߓ��7�%� [�I���Ϧ���o��� �������3�!�W�� ~��G��������� ��	�/�q�V������ w�����������7� .����O�s� ���3�' 79K�o��� ���#//3/5/ G/}/��/�m/�/�/ �/�/??/?�/�/|? �/U?�?�?�?�?�?�? O]?BO�?OuOO�O �O�O�O�O�O5O_YO �OM_;_q___�_�_�_ �__�_1_�_%ooIo 7omo[o}o�o�_�o	o �o�o�o!E3i �o��Y{U�� ���A��h��1� �������������� [�@��	�s�a����� �������3��W�� K�9�o�]��������� ��/�ɯ#��G�5� k�Y���ѯ������ {�����C�1�gϩ� ��ͿW��ϯ������� �	�?߁�fߥ�/ߙ� �߽߫��������Y� >�}��q�_���� ������������� 7�m�[���������� �����!3i W������}�� �/e�� �U����/� /m�d/�=/�/�/ �/�/�/�/?E/*?i/ �/]?�/m?�?�?�?�? �??OA?�?5O#OYO GOiO�O}O�O�?�OO �O_�O1__U_C_e_ �_�O�_�O{_�_�_	o �_-ooQo�_xo�oAo co=o�o�o�o�o) koP�o�q�� ����C(�g� [�I��m�������ُ � �?�ɏ3�!�W�E� {�i�����؟��� ���/��S�A�w��� ��ݟg�ѯc����� +��O���v���?��� ��Ϳ��ݿ��'�i� Nύ�ρ�oϥϓ��� ������A�&�e���Y� G�}�kߡߏ������ �ߵ��߱��U�C�y��g���������$�SERV_MAI�L  ���~��OUTPUT����RV 2�؍�  � (����_���SAVE����TOP10 �2�9� d  	��������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/�}/�/�/�/���YP�|���FZN_CF�G ڍ����j��!GRP� 2��'&� ,�B   A=0��D�;� B>0� � B4��RB{21l�HELL�"C܍�$�L�M�7|�?�;%RSR�? �?�?O�?%OOIO4O mOXOjO�O�O�O�O�O��O_!_3^�  �R3_a_s_AR_� ��{_�R�P)�xWIR2��d�\�]|�Rh6HK 1�v; �_o"ooFo oojo|o�o�o�o�o�o �o�oGBTf~b<OMM �v?��g2FTOV_E�NB��A�$��ROW_REG_UI����IMIOFWD�L�pߥ~@5�WAIT�r�Y�8��r�v@�0�TIM�u7��j�VA��A�>�_UNIT�s��v$�LC�pTRY�w�$���MON_�ALIAS ?e�yH�he��%�7� I�[�i�������� m����
��.�ٟR� d�v�����E���Я� �����*�<�N�`�� q�������̿w��� �&�8��\�nπϒ� ��O���������߻� 4�F�X�j�ߎߠ߲� ���߁�����0�B� ��f�x����Y��� ��������>�P�b� t�������������� (:L��p� ���c��  �6HZl~)� �����/ /2/ D/V//z/�/�/�/[/ �/�/�/
??�/@?R? d?v?�?3?�?�?�?�? �?�?O*O<ONO`OO �O�O�O�OeO�O�O_ _&_�OJ_\_n_�_�_ =_�_�_�_�_�_�_"o 4oFoXooio�o�o�o �ooo�o�o0�o Tfx��G�� ����,�>�P�b� ���������Ώy�����(�:���$S�MON_DEFP�RO ����c� �*SYSTEM�*M�RECALL� ?}c� ( ��}xyzra�te 61=>1�92.168.5�6.1:7188 �� ��Б۟���v�}
��11 �� ��ҟc�u������4� F�X����� ���į ֯g�y�����0�B�T� ���	������ҿc� uχϚ���>�P����� ��*ϼ���_�q߃� �Ϩ�:�L��������߸�360����c��u���tpdiosc 0-�0 ?��Q�������tp?conn 0-ݻ����^�p����0co�py md:pi�ckup.tp �virt:\temp\��0S�������/��lace���0���dv��7���frs:ord�erfil.da�t3mpback@>P����.��b:*.*�0���cu��2x�:1\,�>0 V�(�/�3�a�� :��h/z/�/��: U�/�/
?�/A�/ d?v?�?�,?@/��? �?O/+/�?O/`OrO�O�)� .O@ORO�O��O_��3700 �O�Od_v_�_���� ==<RT_�_�_	o.�_ �_dovo�o�/�/ 6?Ih�o�o�o?$?�o �X�odv��?,�O <RV���O�� >P�h�z����O1�C� U����
��#_��?13924 ԏe�w����c��7�@� R����������Пa�s����g8�o�o�� ?�ۯ���o$��7� ӯd�v����,���:� W����ϟ`4#��� 1�ؿi�{ύϠ���;� V���������B����e�w߉ߚb�$SN�PX_ASG 2��������� >�`%y�����  ?����PARAM ������ �	*��P�d�`��*�����OFT_K�B_CFG  ��c�՞�OPIN_�SIM  ���%������R�VQSTP_DS�Bk�%����SR� �� � }&��ONROD���0���TOP_O�N_ERR  �/�W�L�PTN ����A�H�RING_PR�MV� ��VCNT_GP 2��'��x 	�����``�� ��$��VD��RP 1���(� ��_q��� ����%7 I[m����� ���/!/3/Z/W/ i/{/�/�/�/�/�/�/ �/ ??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_r_o_�_�_�_�_ �_�_�_�_o8o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c����� ������Ϗ���� )�P�M�_�q������� ��˟ݟ���%�7� I�[�m��������ܯ�ٯ����!�3�=P�RG_COUNT�L���[�_�EN�B��Z�M��N䑿_�UPD 1��T  
H��ۿ� ��(�#�5�G�p�k�}� �ϸϳ����� ���� �H�C�U�gߐߋߝ� ���������� ��-� ?�h�c�u����� ��������@�;�M� _��������������� ��%7`[m ������� 83EW�{� �����/// //X/S/e/w/�/�/�/ �/�/�/�/?0?+?=?�O?x?s?�?Q�_IN�FO 1�ɹ�� �F��?�?�?O�9��]MEA?��>>�O�7���PA6�SBʿ�u�P�Y?SDEBUGi�ʰ��0d��z@SP_�PASSi�B?~�KLOG �ɵ+���0>H�?�  ����1U�D1:\�D�>�B_MPC�Mɵ:_L_ɱ��Aj_ ɱVSAV ��MA�A�B��5 XSVnKT�EM_TIME �1��G�� 0*��m��dlXl_�0���T1SVGUNYSİj�'���`�ASK_OPTICONi�ɵ����?a�_DI�@��[eBC�2_GRP 2��ɹ�T�o�1@�  �C��cP��`CFGg �k�\ �V�f`
EOB- Rxc����� ����>�)�b�M� ��q���������ˏ� �(��L�7�p����V n���n�ϟ�\���� �;�&�_�q^�QdT� ������ѯ������ �)�+�=�s�a����� ����߿Ϳ���9� '�]�Kρ�oϑϓϥ� ���Ȭ�����1�C� ��g�U�wߝߋ����� �߳�	���-��Q�?� a�c�u�������� ����'�M�;�q�_� �������������� 7��Oa�� !�����!3 EiW�{�� ���/�///S/ A/w/e/�/�/�/�/�/ �/�/??)?+?=?s? a?�?M�?�?�?�?O �?'OO7O]OKO�O�O �OsO�O�O�O�O_�O !_#_5_k_Y_�_}_�_ �_�_�_�_o�_1oo UoCoyogo�o�o�o�o �o�o�?!?Qc �o�u����� ��)��M�;�q�_� ������ˏ���ݏ� �7�%�G�m�[���� ����ٟǟ����3� !�W�o�������ï A��կ����A�S� e�3���w�����ѿ�� ����+��O�=�s� aϗυϧ��ϻ����� ��9�'�I�K�]ߓ� �߷�m��������#� ��G�5�W�}�k��� ����������1�� A�C�U���y������� ������-Q? uc������ ���/A_q� �����/�� �$TBCSG_GRP 2����  ��  
 ?�  J/\/F/�/j/ �/�/�/�/�/�/;#"�*#�1,d0�?1?!	 HDw 6s33[2g�\5O1B�!�x?�9D)�6L{�ͣ1>���g6Ƙ0CF�?�?�8ff�f�1�>��!OIC�j��6�1H4B�C{OO)HɌ�0|A�]0@HD@O_O)H�1�8CFr�O�M@ �. XU&_�O _Q_n_9_K_�_�_�[�?��0�Sp �	�V3.00�R	�rc65�S	*`�T"o�V|A�0j 8 `�Y G`\mHo  � �%@a�_�o�c#!J2*#��1-�o�hCFG7 ��;!C!�j�B"]b�l|�BPz�P va������ ���<�'�`�K��� o�������ޏɏ�� &��J�5�n�Y�k��� ��ȟ������\	� �-�ן`�K�p����� ����ޯɯ��&�8� �\�G���k�����! /ۿ�����5�#� Y�G�}�kϡϏϱ��� ��������C�1�S� U�gߝߋ��߯����� 	����?�-�c�Q�� ��Y����m������ )��M�;�q�_����� ������������% I[m9��� ����!E3 iW�{���� �/�///?/A/S/ �/w/�/�/�/�/�/�/ ?+?��C?U?g??�? �?�?�?�?�?�?OO 9OKO]OoO-O�O�O�O �O�O�O�O_�O!_G_ 5_k_Y_�_}_�_�_�_ �_�_o�_1ooUoCo yogo�o�o�o�o�o�o �o	+-?uc ����y?��� �;�)�_�M���q��� ����ݏ�����7� %�[�I��������o� ٟǟ����3�!�W� E�{�i���������ï �����A�/�e�S� u����������ѿ� ����+�a��yϋ� ��G��ϻ������'� �K�9�o߁ߓߥ�c� �߷�������#�5�G� ��}�k������ ��������C�1�g� U���y����������� 	��-Q?a� u������� /���q_�� �����/%/7/ �/m/[/�//�/�/ �/�/�/?�/?!?3? i?W?�?{?�?�?�?�? �?O�?/OOSOAOwO eO�O�O�O�O�O�O�O __=_+_M_s_a_�_ C�_�_}_�_�_o 9o'o]oKo�ooo�o�o �o�o�o�o�o# Yk}�I��� ������U�C� y�g���������я�� ��	�?�-�c�Q�s� u��������ϟ�� )�;��_S�e�w�!��� ��˯��ۯݯ�%�� I�[�m��=�����ǿ8���վ  ��� �)���$�TBJOP_GR�P 2�ݵ��  ?���	A�H��O���� ����pXd� ����� � ��,� @��`�	 �D� ��CaDㄈ�`���fff���>��H�ϻ�L{��	�<!a����>���=�B��  Bp��8�C�D�)�U�CQp��D�S�Ι��8y���v� ?������\<���U�n���%�CV+���/���S�D5m�i�{Բ��ع�<����z�>\�>�33C�  �CA��`�K�j���u�bߐ���z�;��9bB�E�>��׵ҳ� C�V���s����&������;��6���%�]�D&� C���������
Ѷ� �?s33����<Z�;u���ff�ҴK������U�)C -_i�u��� ���*Ic M�����Ƙ�����	V3.0}0f�rc65eă* e��/ '� F�  F��� F� F��  G� G�X G'� G;�� GR� Gj�` G�� G��| G� G��� G�8 G��� G�< H�� H� H���2 Ez  E�@ E�� EB �F� FR FZ F��� F� F��P<"G � G�pL#?h GV�� GnH G��� G�� G�(� =u=+U�(�$`Q��?2�3?��  ��M?[:A��*SYSTEM
!�V8.30218� �38/1/20�17 A y � p7M�TP_�THR_TABL�E   $ �$�1ENB��$�DI_NO��${DO�4  ��1�CFG_T � 0�0MAX_I�O_SCAN�2M;IN�2_TI�2D�ME\��0@�0 � � $C�OMMENT w$CVAL	C�T�0PT_IDXꉠEBL�0NUM�QBENDIJfAZIT�ID]B $D�UMMY13���$PS_OVERoFLOW�$�F��0FLA�0YP�E�2�BNC$GLB_TM�7�EF@�1��0ORQCTRL��1�$DEB�UG�CRP�@2@ � $SBR_PAM21_VP� T$SV_E?RR_MODU4S�CL�@RACTI�O�2�0GL_VI�EW�0 4 �$PA$YtRZ�tRWSPtR�A$�CA@A�1"�_SUeU �0N|�P3@$GIF3@}$eQ lP_S�PNiQ LpP�VI<P��PF�RE�VNEA�RPLAN�A$�F	iDISTAN�Cb��JOG_�RADiQ@$�JOINTSP���TMSETiQ�  �WE�UACO�NS2@B�RONF�iQ	� $M�OU1A`�$LO?CK_FOL�A�2oBGLV@CGL�hTEST_XM@@NraEMPE`,R�b<�B`�$US;AfPFH`2P�S�a�b�MP_�`�aQC�ENEdRr $K�ARE�@M�3TP�DRAhP;t2aVEgCLE�32dIU�a�qHE�`TOO�LH`�0qsVI{sR�ESpIS32�y6�4�3ACHX`�`f~qONLE�D29�B��pI�1  @�$RAIL_BO�XEHaPROB�O�d?�QHOW�WAR�0�r�@�qR'OLM�B�A�C ��SK�r�@�0O_F�9�!��S�qiQ
n>o �RVpOCiQ�_�SLOGaK�,�2aQOUZbR�e�AELECTE|<P`�$PIP�f�NODE�r�r�qI�N�q2^��pCOR�DED�`�`}��0P�9P@  D ]�@OBAU`TA �a����C�@���P�q0��ADRA�0F@�TCHup  M,�0EN�2�1A�a�_�Tl�Z@�BObV�WVA!A �� ApeR�5PRE�V_RT�1$E�DIT��VSHWaR9�S@	UАIS`�yQ$IND0@1�QB蓗q$HEA�D�5@ ��p5@��K�EyQ�@CPSPD.�JMP�L�5�0oRACE�4��a�It0S�CH�ANNEzp�	WT'ICK{s�1M`A�0�@�HN�AD0(^�]D�`CG�P���v��0STYf��qLO��A�3B���jP tk 
��Gr�%$���T=PS�!$UNIGa5A�E�0�F�PORT��SQU�5ptR���B�TEsRCJ@*b�TSG� �PP6�$��DE��$`Thq�0OK@>CV�IZ�D�Q�E�APR�AͲ�1旀PU}aݵ_DO�bk�XSV`K�6A�XI��7�qUR_s�E$T�p��*�>�0FREQ_hp<��ET=�P�b�PA�RA`@.P
@�[�N��ATHr�3@�D��s�s�0 �2SR9_Q�0l}��@�1TRQIc��$`�@f��BRup��VE@@^��NOLD��Ap�7a��x@�A��AV_MG�����/����/�D)�D;�DM�J/_ACC.�C��<�9CM��0CYCM@3@��M@_E�����ٺ�@NbSSC�@ o hPDS����1�@SP�0*�AT�:����@��i��BAD�DRES{sB��S�HIF}b�a_2C�H�@&�I�@|��+TV�bI�2]��h�>��C�
�j
�2V8����0 \����A����웱�@��Cn����aºꯆ:R���T�XSCREE�z�0�TINAWS�P;��T�1>�>�jP TQ�7P�B�6Q�P��
��
���RROR_"a�@����E�UEG� �Ⱥ�U��@SXQ�RSyM�� �UNEXg��6��0S_�S�� 	0��>�C�b���o� 26�UE����2GRUͰG�MTN_FLQ��#POHgBBL_r�pWg@�0 ���j�O�Q�LEn����pTO`C�RI;GH�BRDITd��CKGRg@�TE�X,���WIDT�H�sݐB�A�A{q���I_/@H�� � 8 $LT!_ �|�Y0@RyP�b �s�w�B��GOu��0%D0TW� U� �9R�b�LUM�!Ǝ^�ERV��]PFP�`>��1'@r�G�EUR�cF\��Q)&��LP�Z�Ed��)'�$(�$(�p#)U5!+6!+7!+8"�b�>CȰ`��F�qږaS�@EUS=ReT  <��/@qU�R��RFOChq.�PPRIz�m�@?A�� TRIP�qm��UN�0�4!�P` ��0�5��5��b;�5� "T� ̱G �T7���}�&O2OSNAd6RA���;3wq�1#n_�S�^�2H�����aU!"A$�?�?+"��;3OFFT�` P%O��3O@� 1#PD,D$NPGUN#K`S�B_SUBBPk 'SRT�0��&��"a�vp��OR�p�ERA�U���DT�Ib��VsCC��H�' ��C36MFB1����PG?�( (\b`�STE�Qʀ�9PWTѠPE���G�Xd) ����JMOcVE��{Q6RAN4`�?[�3DV�S6RLIM_X�3qV�3qV\XvQ�k\:V1�IP�2V	F��C砽@��G�*��IB�P,�S� _�`�p�b���@/ (0GB�� �"P�@��pr+x# �r �,�tRn�@��s C@TeDRI�PSfQV!�wdԐ���D�$MY_UBY�$\d�;QA�S��q�h�q�bP_S��ף�bL�BMkQ�$j�DEYg�EX�� ���BUM_MUb6�X�D<q US��?��;VGo�PACI�TP�<Uyr�3yr0kSyr:;qREnr�D�1l�8dyr�@,�B/TARGPP�qr8eR{0�@- d�H�;cB	:r��R�D#SWqp�Sn�:s˰�O�!d�Av�3���E���U�p0m��vHK�.��K�AQ���0���?SEA����W�OR�@3��uMRC]Vr/ ��O��M�@C�	ÂC�sÂREF��̆�� gRj�
�� Ȋ�ي�p�=�̆r�_RC�� s�����@����b��8�:bo0 �Т��;��� �e�OU ���r��\c(`+�u���2��<���̰� -�=���f�K�SUL�3a.�C7Po/+p�NT�a��]��a@g��g��!g�&�L�c@���c������!�@)T��s�1���o@�AP_HUR�ۥS]A>SCMP��F�(����_&�R�T������X.��QG�FS�E2d �M� � Y0UF_`�����J��RO� �����W,rUR�GR�mq�I���D_V_h[D�@zY��3�W�IN.rH���X-V@
A�RqR�P�WEw��w�q|c6v,q��RvL�OiPtc�PMc��3ot +=�PA'{ =�CACH6� ���ŵ�,p����K�ۓ�C�QIo�FR"�T8� $֭�$HO�@�R��`�rc��[�֘0p��ڔ�VP�r�����_SZ3p���6����12� ��]p��l�P��WA3�MP�ڮaIMGx���AyD�qIMREٔ^6�_SIZ�P���!po�6vASYNB{UF6vVRTDh��t�F�OLE_2�D�T��t��0C0aU�s��QP�X�ECCU�xVEM�p����#�VIRC��VTP�����G�p��t��LA�s�!��Q�Mco4��;�CKLASQC	��ђ�@�5  �A�� @�&B�T$��$`��6 A|F@o���Xñ�T� o�?a��"�uI���rl/��`BG� VEJ��`PK|p1���֖���HO+��R7 � }F���E�SLOW}w]RO>SACCE*@-�=�xVR:��11�yrcAD�/0rPA�ԩ&�D�1�M_qBa�E��JMP����A8y�b�$SS�C6u��M��C��@9$2��S8��N/�PwLEX��: T��C�Q��6�FLD6?1DEZ�FIQ r�O�qty��BVP2>��;� ϱP�V多�MV_PI Z��G�BP��`а�FIQ�PZ�$��������GA�%p�LOO0Tp�JCBT*����� ��ړPLAN�R&�L��F���cDV�'M �p���U�$�S�P.q �%�!�%#�㱶C4rG����RKE�1�VANC]G�A.0p <�@�?�?R_A�a = �?q??T0�9�)�rG> hܰ�	��K9��fA2b<X@̠OU�e�ݒA��
O���SuK(�M�VIE�p2= S0:�|R�? <{@XMԊ`U�MMY����Re���D��� �@C�U�`b�U�@@ �$�@TIT 1g$PR8�UOPT�VSHIFʀ�A`�a���T��0����$�_R$�UړQ.qZ�U�s �ot�Qav�Q5fS9TG@cVSCO��vQCNT���3� }w�R lW�RzV�R�W�R�XLo�^opjjA2��51D�>a�0� �pS�MO��B%X�J,�@1u���_���@iC%�Gi�LI� ���'��XVR�DD�Y�@T�� ZABCP�E�r�bM��]
��ZIP�EF%���LV��L�����AZMPCF�eG�y�$p?�rDMY_LN$@Ar8��dH ���g���>�MCMİC��COART_Xq�P�1? $JvsptD��|r�r�w���u����UXW�puUXGEUL�x�q�u�t �u�q�q�y�q�v�b�eI Hk�d����Y�`D�� J �8o�	V�EIGH���H?("��f��ĔK �= �C����`$B&�K���1_X�B��LgRV� F^���COVC؀qrfq 9��@}�e�
�����7�D�TRȰ?�V��1�SPH� ǑL� !�S�i�{����S�T�S  �3�����@��@u��<�ѐNa1 ���� ������������������������	���
�����������������;���RDI������ğ֟����t�O|����� ����ίஔ�Sz��� >�����ſ׿��� ��1�C�U�g�yϋ� �ϯ����������v� }���8�!�3�E�W�� �'�9�K�]����[ ����U�5` A;�����0���@A�v�^`BF_TT��ի���I�V>0n�J�_�I�R� 1&� 8�����%к� ��C�  ������������ "�4�F�X�j�|����� ��������1g@BTjx��� ��р����0B QI�ZlJ ��������� /"/4/F/X/FҒ�t/ �/b*���/�/��bv��@`�v�MI_CWHANU� `� #3��dV�`�u�&0ET�>�AD ?��
y0�m��/�/�?�?d�d0RLPs�!&��!�4�?�<SNM�ASKn8��1255.4E0�33OEO�WO�OOLOFS�^Q �`�$X9ORQCTRL &�"V�m��O��T�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo�(l�OKo:ooo��PEΌpTAIL8�JPG�L_CONFIG� 	�ᄀ�/cell/$C�ID$/grp1�so�o�o1�#� �?\n����E ����"�4��X� j�|�������A�S�� ����0�B�яf�x� ��������O����� �,�>�͟ߟt���������ίB�}c��� (�:�L�^���`o��e��b���Ϳ߿��� \�9�K�]�oρϓ�"� �����������#߲� G�Y�k�}ߏߡ�0��� ���������C�U� g�y����>����� ��	��-���Q�c�u� ������:������� );��_q�� ��H��% 7�[m�����]`�User View �i�}}1234567890�
//./�@/R/Z$� �cz/���2�W�/�/�/�/ ??u/�/�3�/d? v?�?�?�?�??�?�.4S?O*O<ONO`OrO�?�O�.5O�O�O�O@__&_�OG_�.6�O �_�_�_�_�_�_9_�_�.7o_4oFoXojo|o�o�_�o�.8#o�o�o�0B�ocir �lCamera��o������NE�,�>� P��j�|�������ď�I  �v�)��&� 8�J�\�n�������� �ڟ����"�4�[��vR9˟�������� ȯگ�����"�m�F� X�j�|�����G�Y�I 7�����"�4�F�� j�|ώ�ٿ�������� ��߳�Y�����Z�l� ~ߐߢߴ�[������� G� �2�D�V�h�z�!� �unY���������� ���B�T�f������ ����������Y�"i{� 0BTfx�1�� ���,> P��Y��i���� ����/,/>/� b/t/�/�/�/�/cu9H/�/?!?3?E?W? �h?�?�?F/�?�?�?��?OO/O�j	�u0 �?jO|O�O�O�O�Ok? �O�O_�?0_B_T_f_ x_�_1OCO�p�{._�_ �_oo+o=o�Oaoso �o�_�o�o�o�o�o �_�u���oOas� ��Po���<� '�9�K�]�o�PEc� ���͏ߏ���� 9�K�]����������� ɟ۟����ϻr�'�9� K�]�o���(�����ɯ �����#�5�G�� ��;�ޯ������ɿۿ ���#�5π�Y�k� }Ϗϡϳ�Z�����J� ���#�5�G�Y� �}� �ߡ������������<���  ��N� `�r���������x����   $� ,�J�\�n��������� ��������"4F Xj|����� ��0BTf x������� //,/>/P/b/t/�/��  
��(  ��B�( 	  �/�/�/�/�/??8? &?H?J?\?�?�?�?�?t�?�*4� �n� O1OCO��gOyO�O�O �O�O��O�O�O_VO 3_E_W_i_{_�_�O�_ �_�__�_oo/oAo So�_wo�o�o�_�o�o �o�o`oroOa s�o������ 8�'�9��]�o��� �������ۏ���F� #�5�G�Y�k�}�ď֏ ��şן�����1� C�U���y�������� ӯ���	��b�?�Q� c�����������Ͽ� (�:��)�;ς�_�q� �ϕϧϹ� ������ H�%�7�I�[�m���� �ߵ���������!� 3�E�ߞ�{����� ����������d�A� S�e������������ ��*�+r�Oa�s������0@ A�������� ��)frh:�\tpgl\ro�bots\r20�00ic6_16?5f.xml�` r�������/����/3/E/W/ i/{/�/�/�/�/�/�/ �//
?/?A?S?e?w? �?�?�?�?�?�?�?? O+O=OOOaOsO�O�O �O�O�O�O�OO_'_ 9_K_]_o_�_�_�_�_ �_�_�__�_#o5oGo Yoko}o�o�o�o�o�o �o o�o1CUg y�������o ��-�?�Q�c�u����������Ϗ���K � 88�?��2�� .�P�R�d��������� �П���(�R�<��^���r�����ܫ�$�TPGL_OUT?PUT ����_ ��� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ������ˠ2345?678901���� ����0�8�����_� q߃ߕߧ߹�Q߽��� ��%�7���}A�i� {����I�[����� ��/�A���O�w��� ������W����� +=����s��� ��e�'9 K�Y����� as�/#/5/G/Y/ �g/�/�/�/�/�/o/ �/??1?C?U?�/�/ �?�?�?�?�?�?}?�? O-O?OQOcO�?qO�O@�O�O�O�OyO֡}��_)_;_M___q_�]@���_�_� ( 	 ���_�_o�_ 5o#oYoGoioko}o�o �o�o�o�o�o/ UCyg���������	�?��Ƭ �-�G�u���c����� ��ߏ���`��,�Ώ P�b�@��������Ο p�ޟ����:�L��� p���$�������ܯ� X���$�Ư�Z�l�J� �����ƿؿz���� �2�DϮ�0�zό�.� ���Ϡ�����b��.� ��R�d�B�tߚ��� ���߄�����<�N� ��r��&������ ��Z�l�&�8���\�n� L����������|��� �� FX��|� 0�����d 0� fxV�� ���//�>/ P/�</�/�/:/�/�/�/�/?
2�$TP�OFF_LIM �[��@W����A2N_SV#0 � �T5:P_M�ON S��74�@�@2�U1S�TRTCHK �S�56_=2VT?COMPATJ8�1�96VWVAR �j=�8N4 R�? O�@}21�_DEFPROG� %�:%CO�NROD�6kO�6_DISPLAY*0��>?BINST_M�SK  �L ~{JINUSER�?΁DLCK�L�KQU?ICKMEN�O�DoSCREPS�~�2tpsc�D��A1P6Y52GP_KYS�T�:59RACE_�CFG �Fr1��4.0	D
?�~�XHNL 2�93��Q�; $B�_�_ o o2oDoVohozj�UITEM 2�[� �%$1234567890�o�e  =<�o�o�os  !{!@�oZC�o{�o� ��9K�o/� �?�e������ #���G���+���O� ��ŏ׏Q�����͟ߟ C��g�y����]��� ���������-���Q� �u�5�G���]�ϯ!� ���ſ)�տ���q� ϕ�����3�ݿ�ϯ� ��%���I�[�m���	� ��c�u��ρ������ 3���W��)��?�� �ߌ��ߧ�����c� S�e�w������k� �������+�=�O��� s�EW��c���� ��9�o ��n����� #�G�"/}=/� M/s/�/��///1/ �/U/?'?9?�/]?�/ �/�/i?�??�?�?Q? �?u?�?PO�?kO�?�O��OO�O)O;O_�TS�R�_UJ�  �bUJ �Q`_UI
 m_�_z_�_8Z�UD1:\�\���QR_GRP �1�k� 	 @`@o!koAo /oeoSo�own��`�o��j�a�_�o�o�e?�  '9{#YG }k������ ���C�1�g�U�w����	�E��ÏSS�CB 2%[ �!�3�E�W�i��{�����\V_CONFIG %]�Q]_�_���OUT?PUT %Y�����S�e�w� ��������ѯ���� �+�_A@�S�e�w��� ������ѿ����� +�<�O�a�sυϗϩ� ����������'�8� K�]�o߁ߓߥ߷��� �������#�5�F�Y� k�}���������� ����1�B�U�g�y� ��������������	 ->�Qcu�� �����) ;L_q���� ���//%/7/H [/m//�/�/�/�/�/ �/�/?!?3?D/W?i? {?�?�?�?�?�?�?�? OO/OAOݟ�>�O �O�O�O�O�O�O�O_ !_3_E_W_J?{_�_�_ �_�_�_�_�_oo/o AoSod_wo�o�o�o�o �o�o�o+=O aro������ ���'�9�K�]�n ��������ɏۏ��� �#�5�G�Y�j�}��� ����şן����� 1�C�U�g�x������� ��ӯ���	��-�?� Q�c�t���������Ͽ ����)�;�M�_� p��ϕϧϹ������� ��%�7�I�[�m�~� �ߣߵ�����������!�3�E�W�i�LH�������s��� hO������1�C�U� g�y���������t��� ��	-?Qcu �������� );M_q�� �����//%/ 7/I/[/m//�/�/�/ �/��/�/?!?3?E? W?i?{?�?�?�?�?�? �/�?OO/OAOSOeO wO�O�O�O�O�O�?�O __+_=_O_a_s_�_ �_�_�_�_�O�_oo 'o9oKo]ooo�o�o�o �o�o�o�_�o#5 GYk}���� ��o���1�C�U� g�y���������ӏ����$TX_SCR�EEN 1������}���&�8�J�\�n��� ������ҟ���� �����P�b�t����� ��!�ίE����(� :�L�ïp�篔����� ʿܿ�e�w�$�6�H� Z�l�~���������� ����� ߗ�D߻�h� zߌߞ߰���9�K��� 
��.�@�R���v��� ����������k����$UALRM_�MSG ?��� ��zJ�\��� �����������������/"SFw+�SEgV  �E���)�ECFG v��  �u�@�  A�  w B��t
 x �s�0BTf�x������G�RP 2� 0�v	 �/+��I_BBL_NO�TE �
T?��l�r���q� +"DEFP�RO5�%9� (%k�/�p�/�/�/�/ �/?�/%??6?[?F?�?j?�?!,INUSER  o-/�?�I_MENHIS�T 18��  �(|  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1`�?`OrO�O�O�)'O~9N381,23�O��O�O	_�O+�O9Ee�ditEBCONRODMOi_{_�__&O>�O138,2�_�_��_o"o�_�_,16�6X_no�o�o�o�@-87oA_SR2,1^o�o 
'o�o;N4]ov�����@'?Q~2 LO�
��.�Q#�0"A �?_�q����������C N������+�=�̏ a�s���������J�ߟ ���'�9�ȟڟo� ��������ɯX���� �#�5�G�֯k�}��� ����ſT�f����� 1�C�U�@�yϋϝϯ� �������	��-�?� Q�c��χߙ߽߫��� ��p���)�;�M�_� q� ���������� ~��%�7�I�[�m��� ���������������� !3EWi{fϟ �����/ ASew��� ���/�+/=/O/ a/s/�/�/&/�/�/�/ �/??�/9?K?]?o? �?�?"?�?�?�?�?�? O#O�?GOYOkO}O�O �O�:O�O�O�O__ 1_4OU_g_y_�_�_�_ >_�_�_�_	oo-o�_ �_couo�o�o�o�oLo �o�o);�o_ q����HZ� ��%�7�I��m���������Ǐ�J�$U�I_PANEDA�TA 1������  �	�}/fr�h/cgtp/w�holedev.stmӏ1�C�U�g�>R�)pri���]�}��Ɵ؟���� � )"�F�-�j�Q� ������į�����ᯀ��B�T�;�x�V����   ��g�����ǿ ٿ����b�3Ϧ�W� i�{ύϟϱ������ �����/�A�(�e�L� �ߛ߂߿ߦ������� ��8���T�Y� k�}�������J� ����1�C�U���y� ��r�����������	 ��-QcJ�n ��0�B��) ;M�q���� ���/h%//I/ 0/m//f/�/�/�/�/ �/�/�/!?3??W?� ��?�?�?�?�?�?:? OO�AOSOeOwO�O �OO�O�O�O�O�O_  _=_O_6_s_Z_�_�_ �_�_�_�_d?v?4O9o Ko]ooo�o�o�_�o*O �o�o�o#5�oY kR�v���� ���1�C�*�g�N� ����o"oӏ���	� �-���Q��ou����� ����ϟ�H���)� �M�_�F���j����� ��ݯį����7��� ��m��������ǿ� ���p�!�3�E�W�i� {�⿟φ����ϼ��� ���/��S�:�w߉��p߭ߔ���D�V�}�����-�?�Q�c�u�) 	��ŉ��������� � ���D�+�h�O�a� �������������� @R9v	�`�Z���$UI_POSTYPE  `��� 	 ����QUICKMEN  ����� REST�ORE 1 `��  �	i�S`N�m~������ /%/7/I/[/�/�/ �/�/�/r�/�/�/j/ 3?E?W?i?{??�?�? �?�?�?�?�?O/OAO SOeO?rO�O�OO�O �O�O__�O=_O_a_ s_�_(_�_�_�_�_�_ �O�_o"o�_Fooo�o �o�o�oZo�o�o�o #�oGYk}�:o ���2���1� C��g�y����������d����	��-��S�CRE� ?��u1scH�u2h�3h�4h�5*h�6h�7h�8h���USERJ�O�a�TLI�j�ksr�є4єU5є6є7є8ё�� NDO_CFG� !����Ѩ P�DATE ����None �_� ��_INFO� 1"`�]�0%3�x�	�f�����˯ ݯ������7��[� m�P�������ǿ�J��OFFSET %�ԿσA֏� *�<�N�{�rτϱϨ� ��Ͼ����A�8� J�w�n߀ߒ������
����UFRA_ME  ʄ��G�RTOL_AB�RT&��>�ENB�G�8�GRP 1&�<Cz  A�����������@������:�� Ug���V�MSK  (j�]�X�N#���]��%�߫��VCCMf�'���RG��E*�	��ʄƉ]D � BH)�p<�2C�)��PN?ـ` ��MR��20���p���"�р	 ����~XC56 �*������N�5р�A@<C�� ��� ʈ);h�c�"�Rр|��Ђ B��� �6�t/T1/ / U/@/y/d/�/�/�/�/ */�/	?�/???�c?\u?��TCC��1��Pf�9�рр��GFS�22w� Й�2345678901�?�2ʈ "�6��?!Oс>,12�$QO_GB@R 8N?:�o=L�� ���������OO A�O�O@O_dOvO�O �O�O�_�O�O�___ �_<_N_`_r_Soeo�_ Ro�o�_�_oo&o8o|��4SELECF��j�$�VIR�TSYNC� ���6�BqSIONT�MOU-tр���cu��3U���U�(�� �FR:\es\+�A�\�o �� �MC�vLOG� �  UD1�vE�X�с' B�@ ����q � ESKTOP-?8U37T7F�6��!�N�`��3�  �=	 1- n6  -��ʆ��xf,p�#�0=�S�ʹ���r�xTRAIN��2�1.��
. d��sq4w (,1��0� �)�;�M�_�q����� ����˟ݟ���I���crSTAT 	5��@�o����E:q$��ۯ�_GE���6w�`. �
���. 2�HOMI�N��7U��U�� �r�a�a�aC�G�um�JMPE�RR 28w
  ʯE:��suTs�� ���߿���'�9�@O�]ώρϓ�_v_�p�RE��9t���LE�X��:wA1-e��VMPHASE'  RuCCb���OFFLpc�<vP2*�t;4�04��8���b@�� �bb>�?s33��Á�1 ��L��ҕԈ�|��t�>x��Â�xf�o.�p��/?P�X� $� 2�x����0� �� �6�+���l��\�j� |���������� � D�V���ZTf��� �������. � ,BPb���� ���//(/:/ �y/�b/��/�/ L/? ??<?n/c?�/ �/�?�?�/�?6?�?�? �?OX?j?\O�?�OJO �?fO�O�O�O�O0O%_ TO_xOm_�O�O�O�_ �_�_�__o>_P_Eo Wo�_xo�_�o�o�o�o���TD_FILTuEt�?�� ��Wp��]o$6HZ l~����� ���)�;�M�_�q�������SHIFTMENU 1@x�<��%����я ��0���f�=�O��� s�����䟻�͟����P�'�	LIV�E/SNAPD�?vsfliv�b����ION �G�U���menu ����:�����±���A���	����b��K��5M����m`@j�����A�pB8�������Ӝѝ������m`� ;ӥ�/�KME��uY��M����MO��B����z��WAITDI/NEND�3����OKN�.�OUT�#��Sa�4�TIM.�����GϮ� @���`ϱ�ϱʞ�2�RELEASE�����TM�����_ACTx��Ȫ��2�_DATA 	C�ի�%i��ߪ����RDIS�b���$XVR2�D���$ZABC_GR�P 1E8�n`,r@h2��ǽZIP1�FD� cCo������x��MPCF_G 1	G8�n`0<o ���=��H8����t� 	|�w�  8R�`����e�����?�k ������5��
\|��  �a  �����7������I��z��YLI�ND�aJ�� ��f ,(  * s�K�p���� �//+.mN/ �r/Y/k/�/��/�/ �/3/?�/�/J?1?n?�U?�/�?�?v�C�2K8��� ��O`o �7O~[Ol�?�Og햨AA�ASPH�ERE 2LS� ?�OX?�O__>_�? �Ot_�_?�_I_/_�_ �_o�_]_:oLo�_�_ �o�_�o�o�o�o#o �$7�ZZ� � k�