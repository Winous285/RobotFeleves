��   ��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A 	  ����PASSNAM�E_T   0� $+ �$'WORD  �? LEVEL � $TI- OU�TT  &F/�� $SET�UPJPROGR�AMJINSTA�LLJY  ?$CURR_O��USER�NUM��STPS_LOkG_P N��$�eT�N�  6 �COUNT_DO�WN�$ENB�_PCMPWD �� DV�IN�!$C� CR=E�PARM:� =T:DIAG:)|�LVCHK!>FULLM0��YXT�CNTD��MENU�A�UTO,�FG_wDSP�RLS��U�fENC/�  CRYwPTE  ����$$CL(   ���;!�� 4D 0 V� IO� :&w+ �
L!�IRTUA� :/��$DCS_COD�@���?%�  {W�'_S  v*%�!x �&�A9�1�"w!� 
 $B!���-�/?  ?6?D?Z?h?~?�?�? �?�?�?�?�?OO2O\,#'SUP� �+04OFO�#FfOxO|�O��  �L��A���O � �� �V�[t&��j���D�ON_���W
_��+!�Ux_UCL�UGH 1w)/ + �)�_ �_�_oo)o;oMo_o qo�o�o�o�'�_�o�o �o/ASew ����o���� �+�=�O�a�s����� ����ߏ���'� 9�K�]�o��������� Ə۟����#�5�G� Y�k�}�������¯ �����1�C�U�g� y���������Я��� 	��-�?�Q�c�uχ� �ϫϽ�̿������ )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{������������� ��/ASew ������%