��  I��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����SBR_T �  | 	$SV�MTR_ID � $ROBOT�9$GRP_�NUM<AXIS�Q6K 6NFF~3 _PARAMF�	$�  �,$MD SPD_[LIT  &2*�� � � � �$$CLAS�S  �������� � � VER�SION��  �
�IRTUAL��' � 1 � T����R-2�000iC/16�5F���  �aiSR22/4�E 80A��
�H1 DSP1-�S1��	P01�.02W,  g	� ��� �  �# ��л��������
�=��r9  �:!a������ @�H+  ����	`� gY�� � ���  }}���������L  2�&����>A�w��u��ψ
"����&���| & ����� �������������+� �����Z�������B� U K ���� �5� :?�����'b�
��c/�/�/�/?��g�?��3<?�a?s?�?��3|2���=f����3x��4+��<����{�Ň����?�?����<N`30/3j2|����ߜ���������~��%����"8 l�� ^�o�������i' � ��&����� 5���:�����A��	���:+��hJ #N ���� ����R�?��}����z'���!�,�c9?	`D 0���� ���#p�"@��x��_�_�_�_�_$3���_B?oo/o  �Z���6<��@����<��g�>3���0�j�cQ�
'�H�o�o�0��?NO�r3|b@OROdK��0tO�O�O�@��G =�'>>�K�4����0���������(:+�  � R__���w���z(��w@_\T_f_x_A�S�e�w�=|���_��я �>o��+�=�O��o��o `10h4�o4|4�o}z�����(�����2�`,8	���� 0��� ��ߍ���b!'6�6�!!p�A�S���- ��/�� l�toc��#����z!��ks��y���c�!�f <�#S ��u�#º'  �
,�����'�9�$3
�>���fd���������ѿ�0���b�t� ��rE5|5����П�U"�����x�����T'#(#�(8�����+�p��z�m�t5�����{�b�� �య%į֯诱�������=���i�2�D� V�h�z������RO@�r6|6dόvψ��P�Ϯ�����	�����'�A�Ϲ���Qd> '	��
P5�M��p#oH�*��4�qq��|ߎߠ�i{��=���/�� 
.@Rdv��?����xTa(��Ng�	�,����/ /2/D/ V/h/z/�/�/�/�/�/��/�/
??.?@?P<� P?t?�?�?�?�?�?�? �?OO(O0C��FO ����O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_o^? &o8oJo\ono�o�o�o �o�o�o6OhOZO#~O �OXj|���� �����0�B�T� f�x�������
o��� ����,�>�P�b�t� �����o����*<N �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�ȏ������ ƿؿ���� �2�D� V�ҟğn������� ����
��.�@�R�d� v߈ߚ߬߾������� ��*N�`�r�� �����������^� �ς�K��ϸπ����� ����������"4 FXj|���� �2��0BT fx������ �R�d�v�>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? ��?�?�?�? OO$O 6OHOZOlO~O���O /"/4/�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRo�? vo�o�o�o�o�o�o�o *�O�O�Os�O �O������� &�8�J�\�n������� ��ȏڏ���Zo�4� F�X�j�|�������ğ ֟�D� �z�� f�x���������ү� ����,�>�P�b�t� ������������ �(�:�L�^�pςϔ� ��"����8�J�\�$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�ֿ������� ����
��.�@�R��� ���ϛ���������� *<N`r� ������ &��8\n��� �����/l�5/ (/�������/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? @OO,O>OPObOtO �O�O�O�O�OJ/</�O `/r/�/L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�? �o�o�o�o 2D Vhz�O_�O�_ 0_�
��.�@�R�d� v���������Џ�� ��*�<�N��o`��� ������̟ޟ��� &�8��]�P���� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ����h�0�B�T� f�xϊϜϮ������� ��r�d�߈�����t� �ߘߪ߼�������� �(�:�L�^�p��� �����&��� ��$� 6�H�Z�l�~������� 0�"���F�X� 2D Vhz����� ��
.@Rd v������� //*/</N/`/���/ x/���/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O �XOjO|O�O�O�O�O �O�O�O__�/�/6_ �/�/�/�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�oNO (:L^p�� ���&_X_J_�n_ �_H�Z�l�~������� Ə؏���� �2�D� V�h�z������o��ԟ ���
��.�@�R�d� v���������,�>� ��*�<�N�`�r��� ������̿޿��� &�8�J�\ϸ��ϒϤ� �����������"�4� F�¯��^�د����� ��������0�B�T� f�x���������� ����v�>�P�b�t� ��������������N� ��r�;�ߨ�p�� ����� $ 6HZl~��� �"���/ /2/D/ V/h/z/�/�/�/�/ �/BTf.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O ��O�O�O�O�O__ &_8_J_\_n_�/�/�_  ??$?�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0B�O fx������ ���v_�_�_c��_ �_������Ώ���� �(�:�L�^�p����� ����ʟܟ�J �$� 6�H�Z�l�~������� Ưد4����j�|��� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬ�������� ��*�<�N�`�r߄� ������(�:�L�� &�8�J�\�n���� �����������"�4� F�X�j��ώ������� ������0B�� ���ߋ������� �,>Pbt �������/ /r�(/L/^/p/�/�/ �/�/�/�/�/ ?\%? ?���~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O 0/�O
__._@_R_d_ v_�_�_�_�_:?,?�_ P?b?t?<oNo`oro�o �o�o�o�o�o�o &8J\n���O ������"�4� F�X�j��_�_�_��o  o�����0�B�T� f�x���������ҟ� ����,�>��P�t� ��������ί��� �(���M�@���̏ޏ ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������X� �2�D� V�h�zߌߞ߰����� ��b�T���x�����d� v����������� ��*�<�N�`�r��� ����������� &8J\n����  ���6�H�"4 FXj|���� ���//0/B/T/ f/��x/�/�/�/�/�/ �/??,?>?P?�u? h?���?�?�?O O(O:OLO^OpO�O�O �O�O�O�O�O __$_ �/H_Z_l_~_�_�_�_ �_�_�_�_o�?|?&o �?�?�?�o�o�o�o�o �o�o
.@Rd v������>_ ��*�<�N�`�r��� ������oHo:o�^o po8�J�\�n������� ��ȟڟ����"�4� F�X�j�|������į ֯�����0�B�T� f�x�ԏ����
��.� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�Lߨ�p߂ߔ� �߸������� ��$� 6ﲿ��N�ȿڿ쿴� ��������� �2�D� V�h�z����������� ����
f�.@Rd v������>� p�b�+���`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/?"?4? F?X?j?|?�?�?��? �?2DVO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �/�_�_�_�_�_�_o o(o:oLo^o�?�?vo �?OO�o�o $ 6HZl~��� ����� �2��_ V�h�z�������ԏ ���
�fo�o�oS��o �o��������П��� ��*�<�N�`�r��� ������̯ޯ:��� &�8�J�\�n������� ��ȿ$���Z�l�~� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ��������� ����,�>�P�b�t� ��������*�<�� �(�:�L�^�p����� ���������� $ 6HZ��~��� ���� 2�� ���{������ ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ?b?<?N?`?r?�? �?�?�?�?�?�?LO O���nO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_  ?�_�_oo0oBoTo foxo�o�o�o*OO�o @OROdO,>Pbt �������� �(�:�L�^�p����_ ����ʏ܏� ��$� 6�H�Z��o�o�o���o ؟���� �2�D� V�h�z�������¯ԯ ���
��.���@�d� v���������п��� ��t�=�0Ϫ���Ο �ϨϺ��������� &�8�J�\�n߀ߒߤ� ��������H��"�4� F�X�j�|������ ��R�D���h�zό�T� f�x������������� ��,>Pbt ������� (:L^p��� ���&�8� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?�h?�?�?�?�?�? �?�?
OO.O@O�eO XO����O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo p?8oJo\ono�o�o�o �o�o�o�o�ozOlO �O�O�O|���� �����0�B�T� f�x���������ҏ.o ����,�>�P�b�t� ������8*�N `(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~�ڏ���� ƿؿ���� �2�D� V�h�ğ�π����� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<`�r�� ������������ &��ϔ�>������Ϥ� ����������"4 FXj|���� ���V�0BT fx�����.� `�R�/v���P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�? OO$O 6OHOZOlO~O�O��O �O"/4/F/_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo �?�o�o�o�o�o�o�o *<N�O�Of �O�O_����� &�8�J�\�n������� ��ȏڏ����"�~o F�X�j�|�������ğ ֟���V�zC�� �x���������ү� ����,�>�P�b�t� ��������ο*��� �(�:�L�^�pςϔ� �ϸ������J�\�n� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z��述����� ����
��.�@�R�d� v����ώ���,��� *<N`r� ������ &8J��n��� �����/"/~� ����k/�����/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?RO,O>OPObOtO �O�O�O�O�O�O</_ �Or/�/�/^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o O�o�o�o 2D Vhz��__� 0_B_T_�.�@�R�d� v���������Џ�� ��*�<�N�`�r��o ������̟ޟ��� &�8�J�������  �ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����z�0�T� f�xϊϜϮ������� ���d�-� ߚ����� �ߘߪ߼�������� �(�:�L�^�p��� �������8� ��$� 6�H�Z�l�~������� ��B�4���X�j�|�D Vhz����� ��
.@Rd v������� //*/</N/`/r/��  ���/(�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FO�XO|O�O�O�O�O �O�O�O__0_�/U_ H_�/�/�/�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o `O(:L^p�� �����j_\_� �_�_�_l�~������� Ə؏���� �2�D� V�h�z������� ���
��.�@�R�d� v������(���>� P��*�<�N�`�r��� ������̿޿��� &�8�J�\�n�ʟ�Ϥ� �����������"�4� F�Xߴ�}�p����� ��������0�B�T� f�x���������� ����,���P�b�t� �������������� �߄�.�ߺ��ߔ ����� $ 6HZl~��� ���F�/ /2/D/ V/h/z/�/�/�/�/ PB?fx@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O��O�O�O�O__�&_8_J_\_n_�_�%��$SBR2 1� 5�P T0? � �C?7 �_�_�_o o2oDo Vohozo�o�o�o�o�o�Q�o�_!3E Wi{����� ���o� A�S�e� w���������я��� ��+��O�2�s��� ������͟ߟ��� '�9�K�]�@���d��� ��ɯۯ����#�5� G�Y�k�}���r����� ׿�����1�C�Uπg�yϋϝϯ��Ϥ�~ �_�����!�3�E�W� i�{ߍߟ߱������� �����(�:�L�^�p� ����������� � ����H�Z�l�~��� ������������  2D(�:�z��� ����
.@ RdvZ���� ��//*/</N/`/ r/�/�/�/��/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�/�?O "O4OFOXOjO|O�O�O �O�O�O�O�O_�?0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>o"_ boto�o�o�o�o�o�o �o(:L^p To������ � �$�6�H�Z�l�~��� ���Ə؏���� � 2�D�V�h�z������� ������
��.�@� R�d�v���������Я ���؟�*�<�N�`� r���������̿޿� ��&�
�4�\�nπ� �Ϥ϶���������� "�4�F�X�<�|ߎߠ� ������������0� B�T�f�x��n߮��� ��������,�>�P� b�t������������� ��(:L^p ��������� $6HZl~� ������/ / D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?6/v?�?�?�?�?�? �?�?OO*O<ONO`O rOV?h?�O�O�O�O�O __&_8_J_\_n_�_ �_�_�O�O�_�_�_o "o4oFoXojo|o�o�o �o�o�o�_�o0 BTfx���� �����o,�>�P� b�t���������Ώ�� ���(�:��^�p� ��������ʟܟ� � �$�6�H�Z�l�P��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ���&�8�J�\�n�� ������������� "���X�j�|����� ����������0 BT8�J����� ���,>P bt�j���� �//(/:/L/^/p/ �/�/�/�/��/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�/O O 2ODOVOhOzO�O�O�O �O�O�O�O
__ O@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo2_ ro�o�o�o�o�o�o�o &8J\n� do������� "�4�F�X�j�|����� ���֏�����0� B�T�f�x��������� ҟ��ȏ��,�>�P� b�t���������ί� �����:�L�^�p� ��������ʿܿ� � �$�6��D�l�~ϐ� �ϴ���������� � 2�D�V�h�Lόߞ߰� ��������
��.�@� R�d�v���~߾��� ������*�<�N�`� r��������������� &8J\n� ��������� "4FXj|�� �����//0/ T/f/x/�/�/�/�/ �/�/�/??,?>?P? b?F/�?�?�?�?�?�? �?OO(O:OLO^OpO �Of?x?�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�O�O�_�_o o 2oDoVohozo�o�o�o �o�o�o�_�o.@ Rdv����� �����o<�N�`� r���������̏ޏ�� ��&�8�J�.�n��� ������ȟڟ���� "�4�F�X�j�|�`��� ��į֯�����0� B�T�f�x��������� ҿ�����,�>�P� b�tφϘϪϼ����� Ŀ��(�:�L�^�p� �ߔߦ߸������� � ���6�H�Z�l�~�� ������������ � 2��(�h�z������� ��������
.@ RdH�Z����� ��*<N` r��z���� //&/8/J/\/n/�/ �/�/�/�/��/�/? "?4?F?X?j?|?�?�? �?�?�?�?�?�/O0O BOTOfOxO�O�O�O�O �O�O�O__,_OP_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^oB_ �o�o�o�o�o�o�o  $6HZl~� to������ � 2�D�V�h�z������� ����
��.�@� R�d�v���������П �Ə؏�*�<�N�`� r���������̯ޯ� ����
�J�\�n��� ������ȿڿ���� "�4�F�*�T�|ώϠ� ������������0� B�T�f�x�\Ϝ߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� �������� 2DVhz��� ����
//./@/ $d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?V/�?�?�?�?�?�? OO&O8OJO\OnO�O �Ov?�?�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�O�O�_oo0o BoTofoxo�o�o�o�o �o�o�o�_,>P bt������ ���(�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�