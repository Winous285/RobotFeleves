��   b�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����CELLSET�_T   �w$GI_STY�SEL_P }7T  7ISO:iRibDiTRA�R�>�I_INI; �����bU9AR�TaRSRPNS�1Q234�5678�Q
TROBQACKSNO� �)�7�E�S �a�o�zU2 3 4 5 6 7 8awn&GINm'D�&��) %��)4%��)P%�̖)l%SN�{(OU���!7� OPTNAA�73�73.:B<;�}a6.:C<;CK;C�aI_DECSN�A�3R�3�TRY�1��4��4�PTHCN�8D�D�INCYC@HG��KD�TASKOK �{D�{D�7:�E� U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V�8�Tb@SEGq�Tp��T�@REQ� d�drG�:Mf�GJO_HFAUL�Xpd�dvgALE�  �g�c�g�cvgE� �H<�dvgNDBR�H�dgRGAB�Xtb�p�CLML�Iy@   �$TYPESI�NDEXS�$$�CLASS  O���lq�����apVERSIO�Nix  ��
}qIRTU�ALi{q'61�r���p��q�t+ �UP0 �x�Style Se�lect 	  ����r�uReq. _/Echo����Ack���I?nitiat�p�r��
�^�m�������	��
��  U�������������χ�q)���Option b�it A<��p�B���C4�Deci�s�codY��Tryout mj��6�Path se}gh�ntin.8��Ig�ycX�:�Ta�sk OK��?�M�anual op�t.r�A���B����C� dec�sn ��$�Rob�ot inter�lo7�@�\� isSolQ�4�C��iM�<@���ment<�)��������Ě}�sta�tus=�	MH ?Fault:����Aler�1�C��pn@r 1�z j��;�y���I�; LE_�COMNT ?>�y�   Չ� ѿ�����*�<�N� `�rυϖϨϺ����� ����&�9�J�\�n� �ߒߤ߶����������"�����U��Ђ���Ŵ   ��ENA/B  ��:�����������ꮵM�ENU\��y��NA�ME ?%��(%$*R�זb��P��� t��������������� +O:s^p� �����  $6HZ�~�� �����/ /Y/ D/}/h/�/�/�/�/�/ �/�/?
?C?.?@?R? d?v?�?�?�?�?�?�? �?OM