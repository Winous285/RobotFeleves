��   u��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����UI_CONF�IG_T  �� A$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]2�ODE�
3CWFOCA �4C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"��%�!BA�!j ?Ɵ"BG�%�!jIN=SR$IO}7�PM�X_PKT��"IHELP� M{ER�BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�; } &USTOM0� t $} R?T_SPID�,D�C4D*PAG� ?�^DEVICE�PISCREuEF���IGN�@$FLAG�@C�1 � h 	$PWD_ACCES� E �8��C�!~�%)$LABE� O$Tz j�@��3�B�	CUSR�VI 1  < �`�B*�B��APRI�m� t1RP�TRIP�"m�$�$CLA�@ ����sQ��R��R�hP\ SI�qW  �
�QIRTs1q_�P'2 �L3hL3!p�R	_ ,��?2����Q�P�R�T��Q�R���P�  �T/o��
 ��zQQocouo�o�o�o�o Mo�o�o *<�o`r�� ��I����&� 8�J��n��������� ȏW�����"�4�F� Տj�|�������ğ֟ e�����0�B�T�� x���������үa������,�>�P�b��P�TPTX��p򨅿���P sm����$/soft�part/gen�link?hel�p=/md/tpmenu.dgd� ���"�4��X�j�|� �Ϡϲ�A�������� �0߿�A�f�xߊߜ� ����O�������,�,>����zQ'`V�8	bbS� ($�ߕ�@����������zQ@�Q�c������*k
m�d���
e@� ��P����D@�*dn���	b�#`  �V�������SB 1�XR/ \ }%`�REG VE�D�� who�lemod.ht}m4	singlE�doub\�triptbrows�@�!� ���/AS�|�/Adev�.sJl�o�1�	t���w� G/Y/k/5/�/�/�/�/�/ ?� �P?*? <?N?`?r?�?�?�?�? �6�@?�?�?�? O2O DOE	�/�/wO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ ��_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o	-??z �������
� �O@�R�!�3����� QOcOI�ݏ��*� %�7�I�r�m������ ��ǟٟ�����_/� )�W�i�{�������ï կ�����/�A�S� e�w�����iֿ��� ��0�B�T�f�x�s� �Ϯ�}Ϗ����ϭ��� ��>�9�K�]߆߁ߓ� ������������#� 5�^�Y�k�9����� ����������1�C� U�g�y����������� ����ſ2DVhz ��������
 ��@R	��� ������/*/ %/7/I/r/m//�/�/ �/�/���/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO !�O�O�O�O�O�O�O __0_+T_f_5_G_��_�_�Z�$UI_�TOPMENU �1�P�Q?R 
d�QfA�)*defau�ltqOZM*level0 *\K�	 o� So��_Qocbtpio[�23]�(tpst[1�heo�ouo3o�Eo�-
h58E0�1.gif�(	menu5&ypHqC13&zGr%zEt4M{4�a������ ���eB�C�U�g��y�����,�pri�m=Hqpage,?1422,1��ݏ ���%�0�I�[�m�������2���class,5�������)�4���13�0�f�x�������5���53ʏ���� �2�5���8ٯm�� ������4�ٿ����!�3�^I�P�Q�_kπm]��a[ϕ�o�ft�y�m�o�amf[0��o��	��c[164�g.�59�h�a�L��tC8$|Gr2u K}��azmWw%{�ߩs K�]�6�H�Z�l�~�ɿ ����������𢡊��80$�?�Q�c�u�����̐2���������� 	��ʟ?Qcu� (T�������Ѥ1.�N`r�������ainedic����//���config�=single&>��wintpĀ / `/r/�/�/]J�QV¤/ �/e�/�o�o??1? D?U?g?y?�?�/�?�? �?�?�?	OO-O?O� aO�O�O�O�O�O�O�� __*_<_N_`_�O�_ �_�_�_�_�_m_�_o &o8oJo\ono�_�o�o �o�o�o�o{o"4 FXj�o|��� �����0�B�T� f�x��������ҏ���MNS�,�wω¯����w���s��<�����ϡ�u�͔�V�|�F7��7����԰�Οp�4�ߔ�6��u7���  �����/�A��227쯃�������˿ Z�l�����,�>�P�
/!$13�ϛϭ� ���ϐ�����+�=� O���s߅ߗߩ߻��� ��"���'�9�K�]�����6d��������,$۬74r��/��A�S�e��,����%	�TPTX[209�����24����������18�������(
����0P2���10_��E�tv������Q�u10�1�=�ïqC:4$tre�eviewA#�3��&dual=o�U81,26,4 ����n���� 	//-/�Q/c/u/�/H�/�/ֺ;@b�3` r�?)?;?F/_?q?��?�?�?�?�/�/\2�/t2��O1OCO�?��1�/E���O�O�O�6XO��edit �zO�O_._@_׹? ���OCL_�_�_�_~� �_�_G�o}o�Co Uogoyo�o�o�o�o/o �o�o	-?Qd uӥ������ �I?2�D�V�h�z��� ���ԏ���
��� �@�R�d�v�����)� ��П�������<� N�`�r�����%���̯ ޯ���&���J�\� n�������3�ȿڿ� ���"��_�_X�o|� �o��ϱ��������� �ߋ�)�S�e�x߉� �߭߿��ߓ��,� >�P�b�t￿���� ��������(�:�L� ^�p������������ �� ��$6HZl ~������ � 2DVhz� �����
/� ./@/R/d/v/�/7�I� �/m��/I���??)? ;?M?`?q?�?�/�?�? �?�?�?OO%O7O�� nO�O�O�O�O�O�O%/ �O_"_4_F_X_�O|_ �_�_�_�_�_e_�_o o0oBoTofo�_�o�o �o�o�o�oso, >Pb�o���� �����(�:�L� ^�p��������ʏ܏ /�/$��/H��?MO k�}�������ş؟� W����1�C�U�h�y� ����_Oԯ���
�� .�y�@�d�v������� ��M������*�<� ˿`�rτϖϨϺ�I� ������&�8�J��� n߀ߒߤ߶���W��� ���"�4�F���X�|� ��������e������0�B�T���*defaulta��2�*level�8���������{� �tpst[1�]��ytpio[23���u������	m�enu7.gif��
�13�	�5��
��
�4�u6 �
ʯ?Qcu�� �����//� ;/M/_/q/�/�/�/6"�prim=�p�age,74,1��/�/�/??+?6"��&class,130?f?x?�?�?�?=?O25�?�?�?O O2O5#D<�?lO~O�O�O�O�/�"18�/�O_ _'_9_DON26@_u_��_�_�_�_��$U�I_USERVI�EW 1���R 
����_>��_
o�m (oQocouo�o�o<o�o �o�o�o�o);M _qo~��� ���%��I�[�m� �����F�Ǐُ��� ���.�@���{��� ����ßf������ /�ҟS�e�w�����F� P���̯>���+�=� O�a����������Ϳ p����'�9��F� X�j�ܿ�Ϸ������� ���#�5�G�Y�k�� �ߡ߳����߂����� �z�C�U�g�y��.� ������������-� ?�Q�c�������� ������)��M _q��8��� ��� 2�m ���X��� /!/3/�W/i/{/�/ �/J�/�/�/B/?? /?A?S?�/w?�?�?�? �?b?�?�?OO+O�/ �?JO\O�?�O�O�O�O �O�O�O_'_9_K_]_  _�_�_�_�_�_lX