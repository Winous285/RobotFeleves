��   �A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ��
��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP���HOv��NT. 4� �H�9ADDRT�YP� A H� NG#THOG��z +�LS/ D $ROBOTIG �BPEER�� MwASK@MRU~;OMGDEVK%�RCM+�� :$�� ��QwSIZNTIM�$STATUS�_�?MAILS�ERV�  $PL�ANT� <$LI}N�<$CLU���f<$TOcP$�CC5&FR5&J�EC!�ENB{ � ALAR��B�TP�w#�V�8 S��$VAR)M�ONt&��t&oAPPLt&PA� 8u%�s'POR ��_T!["ALERT�5&2URL }}�#ATTAC[�0ERR_THRO�#US29�38� �CH- �[4MAX�?WS_1�Ny1MOD�z1I� �$y2 � (y1PoWD  ; LAu�00�NDq1TRY�6DELA�3z0�>�1ERSIS�!�2v�RO�9CLK�8qM� ��0XML+ ��#SGFRM�#T�CP�OU�#PI�NG_RE�5OP �!UF�#[A�C�"u%_B_AUZ�@��B~�!DUMMY1�j�A2?>�DM*}� $DIS��� �SM�� l5�!,"%,�'NICCb%H � �0VR#01UP*_D�LVPAR���J@Io/ 3 $�ARP�)_IP�FOW_��F7_INFAD� ܛHO_� IN{FO��TELsG	 P~����� WOR�1$A7CCE� LV�[:�"�ICE�0 a�  �$�S  ����@a��
���
5`PSlA>g  �PbI0AL=oOa'0 V^h
���F����i`�b�e��� ęm��!Ga�o���$�ETH_FLTRs  ]i�` ��������{�� ��m2{�RSHcPD� 1�i  P�o��d��� ����:��F�!� o���W���{�܏�� � Ï$����Z��~�A� ��e�Ɵ�������� � �D��h�+�a����� ¯��毩�
�ͯ�� ?�d�'���K���o�п ������ɿ*��N�� r�5ϖ�Y�k��Ϗ��� �����8���1�n�]�`��U߶�wz _L�1�1}x!1."��0��y���1�y�255.9�����ܶe��2���m� �.�@�R�d�3n��@��������d�4���]���0�B�d�5 ^��������������6���M �� 2�����6AMY�� MY����p{�K`� 'Q� ��~<� /SewJ��v�P���/�%/ 7/I/[///�/�/~t/uٹe�/�,�/i/�2?D?V?h?}�}i�RConnect�: irc�4//?alertsm?�? �?�?�?x5,?O#O5OPGOYOkO}��cd�`pd��pO�O�O�O �O�O __$_6_H_Z_�l_~_{�$ O�_`p( �_�_$?�_oo+oy�):`p���\b��jNeKabe|�Su� D�M�c�n�$SM&Iu�{��%�_�o�$`p�o}��o8�#\�,��TCPIP�b�m�(�~q�EL��	�eSa�  H!TPh�s�rj3_t�p�Bp|��Pq!KCL��{P��>f!CRT@�.������!CON�S���z�qsmo	n���