��   �A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ��
��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP� HOv��NT. 4� �H�9ADDRT�YP� A H� NG#THOG��z +�LS/ D $ROBOTIG �BPEER�� MwASK@MRU~;OMGDEVK����RCM+� :$�� ���QSIZNTIM�$STATU�S_�?MAIL�SERV�  $P�LANT� <$L�IN�<$CLU���f<$TOcP7$CC5&FR5&�JEC!�EN�B � ALAR�B�TP�w#��V8 S��$VA5R)M�ONt&���t&APPLt&PAp� u%�s'POR ��_T!["ALER�T5&2URL �}�#ATTAC�[0ERR_THRO�#US29�38ƚ CH- �[4MA�X?WS_1��y1MOD�z1IF� $y2 � (y1�PWD  ; LA�u00�NDq1TR=Y�6DELA�3z0|��1ERSIS�!�2�RO�9CLK��8M� ��0XML|+ �#SGFRM�#�TCP�OU�#P�ING_RE�5OAP�!UF�#[A�C�"u%_B_AUZ�@���B�!DUMMY1԰�A2?�DM�*� $DISL��SM�$l5��!,"%�'NICC"b%H � 0VR#01U�P*_DLVP+AR��J@Io/ }3 $ARP��)_IPFOW_x��F_IN�FAD� �HO�_� INFO��wTELs	 P~���� WOR~�1$ACCE� �LV�[�"�IcCE�0 a���$�S  ���@aJ��
��
5`PSlA�>g  5�PbI0AL=oOaX'0 ^h
���F��a��i`�b�e��� �m��!Ga�o����$ETH_FL�TR  ]i�` Z�@ % ����{��� �m2{�RSH�cPD 1�i G P�o��d� ������:�� F�!�o���W���{�܏ �� �Ï$����Z�� ~�A���e�Ɵ������ �� ��D��h�+�a� ����¯��毩�
�ͯ ��?�d�'���K��� o�п������ɿ*�� N��r�5ϖ�Y�k��� ���ϳ����8���1߀n�]ߒ�U߶�wz _�L�11}x!�1.��0��y���1|�y�255.9�L����ܶe��2�߀�m��.�@�R�d�3 n����������d�4���]���0�B�d�5^��������������6���M ��� 2����6A�MY� MY����p{�K`�� Q� ��~< �/SewJ��v�P���/ �%/7/I/[///�/�/~t/uٹe�/�,��/i/2?D?V?h?}�}�iRConnect: irc�4�//alerts m?�?�?�?�?x5,?O@#O5OGOYOkO}��c9d�`pd��pO�O �O�O�O�O __$_6_ H_Z_l_~_{�$ O�_`p(�_�_$?�_oo�+oy�:`p�� �\b�jNeKabe|�Suֿ DM�c�n�$�SMIu�{��%�_�o�$`p�o}���o8#\�,��TCWPIP�b�m�(,�~qEL��	�eSa��  H!T�Phs�rj3�_tp�Bp|��Pq!KCL��{P|��>f!CRT@��.�����!C�ONS���z�qs'mon���