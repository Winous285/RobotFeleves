��   �A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ��
��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP� HOv��NT. 4� �H�9ADDRT�YP� A H� NG#THOG��z +�LS/ D $ROBOTIG �BPEER�� MwASK@MRU~�OMGDEVK"� RCM+� :$�� ���QSIZNTIM�$STATU�S_�?MAIL�SERV�  $P�LANT� <$L�IN�<$CLU���f<$TOcP7$CC5&FR5&�JEC!�EN�B � ALAR�B�TP�w#��V8 S��$VA5R)M�ONt&���t&APPLt&PAp� u%�s'POR ��_T!["ALER�T5&2URL �}�#ATTAC�[0ERR_THRO�#US29�38ƚ CH- �[4MA�X?WS_1��y1MOD�z1IF� $y2 � (y1�PWD  ; LA�u00�NDq1TR=Y�6DELA�3z0|��1ERSIS�!�2�RO�9CLK��8M� ��0XML|+ �#SGFRM�#�TCP�OU�#P�ING_RE�5OAP�!UF�#[A�C�"u%_B_AUZ�@���B�!DUMMY1԰�A2?�DM�*� $DIS���� SM�C l5�!,"%�'NICCb%H � 0V�R#01UP*_DLVPARN� J@�Io/ 3 $A�RP�)_IPF�OW_��F_INFAD� ��HO_� INF�O��TELs	# P~���� �WOR�1$ACCE� LV�[�"�ICE�0 a����$�S  �S��@a��
��
5`�PSlA>g�  �PbI0A�L=oOa'0 ^h
�
��F����i`�b�e���� �m��!�Ga�o���$ETH_FLTR  ]iΤ` ���@ �B���{�� �m2{��RSHcPD 1>�i  P�o��d������ �:��F�!�o���W� ��{�܏�� �Ï$�� ��Z��~�A���e�Ɵ �������� ��D�� h�+�a�����¯��� ��
�ͯ��?�d�'� ��K���o�п������ ɿ*��N��r�5ϖ� Y�k��Ϗ��ϳ���� 8���1�n�]ߒ�U߶�lwz _L�11}_x!1.��0���y���1�y�25c5.9�����ܶe��2���m��.�@�R�d�3n�����������d�4���]���0�B�d�5^���� ����������6���@M �� 2�����6AMY� M?Y���p{��K`� Q� ��~<�/S@ewJ��v�P� ��/�%/7/I/[/ //�/�/~t/u� �e�/�,�/i/2?D?V?�h?}�}iRCo�nnect: i�rc�4//alertsm?�?�?�?�? x5,?O#O5OGOYOkO�}��cd�`pd��pO�O�O�O�O�O _ _$_6_H_Z_l_~_{�$ O�_`p(�_�_$? �_oo+oy�:`p���\b�jNeKa�be|�Su� DM�c��n�$SMIu��{��%�_�o�$`p �o}��o8#\�,���TCPIP�bb�m�(�~qEL���	�eSa�  H�!TPhs�?rj3_tp�Bp|���Pq!KCL���{P��>f!C�RT@�.�����?!CONS���z=�qsmon���