��   �A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ��
��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP� HOv��NT. 4� �H�9ADDRT�YP� A H� NG#THOG��z +�LS/ D $ROBOTIG �BPEER�� MwASK@MRU~�OMGDEVK� RCM+� :$�� ���QSIZNTIM�$STATU�S_�?MAIL�SERV�  $P�LANT� <$L�IN�<$CLU���f<$TOcP7$CC5&FR5&�JEC!�EN�B � ALAR�B�TP�w#��V8 S��$VA5R)M�ONt&���t&APPLt&PAp� u%�s'POR ��_T!["ALER�T5&2URL �}�#ATTAC�[0ERR_THRO�#US29�38ƚ CH- �[4MA�X?WS_1��y1MOD�z1IF� $y2 � (y1�PWD  ; LA�u00�NDq1TR=Y�6DELA�3z0|��1ERSIS�!�2�RO�9CLK��8M� ��0XML|+ �#SGFRM�#�TCP�OU�#P�ING_RE�5OAP�!UF�#[A�C�"u%_B_AUZ�@���B�!DUMMY1԰�A2?	�DM�*� $DIS�����SM�C l5�!,"%�'NICCb%H � 0V�R#01UP*_DL�VPARN��J@Io/ 3 �$ARP�)_IPFOW_��oF_INFAD�� �HO_� I�NFO��TEL�s	 P~��܊� WOR�1$oACCE� LV�t[�"�ICE�0� a �$�S ? ���@a��%
��
5`PSlA>g�  �PbI0AL=oOa'�0 ^h
���F��0��i`�b�e���� �m��!Ga�o����$ETH_FLTgR  ]i�` �+ ������{�d� �m2{�RSHcP�D 1�i # P�o��d�� �����:��F� !�o���W���{�܏��  �Ï$����Z��~� A���e�Ɵ��������  ��D��h�+�a��� ��¯��毩�
�ͯ� �?�d�'���K���o� п������ɿ*��N� �r�5ϖ�Y�k��Ϗ� �ϳ����8���1�n��]ߒ�U߶�wz _L��11}x!1E.��0��y���1�>y�255.9���&��ܶe��2���@m��.�@�R�d�3n����������d�4 ���]���0�B�d�5^��������������6���M �� �2����6AM�Y� MY����p{�K`� OQ� ��~<� /SewJ��v�P���/� %/7/I/[///�/�/~t/uٹe�/�,�/�i/2?D?V?h?}�}�iRConnec�t: irc�4//alertsm? �?�?�?�?x5,?O#O�5OGOYOkO}��cd�`pd��pO�O�O �O�O�O __$_6_H_Z_l_~_{�$ O�_`p(�_�_$?�_oo+oRy�:`p��� \b�jNeKabe|�Su� �DM�c�n�$SMMIu�{��%�_�o�$`p�o}��o�8#\�,��TCP+IP�b�m�(��~qEL��	�eSa��  H!TP�hs�rj3_�tp�Bp|��Pq!KCL��{P��>>f!CRT@�.������!CO�NS���z�qsmon���