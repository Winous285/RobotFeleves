��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�   � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d PPINFwOEQ/ ��L A �!�%/� H� �&�)EQUIP 2� �NAMr �'2_�OVR�$VEgRSI3 �� COUPLED�w $!PP_� OCES0s!_81s!͗!PC> �!� � $SOF�T�T_IDk2TOTAL_EQs 3$�0�0NO�2U �SPI_INDE�]�5Xk2SCRE�EN_(4_2SI�GE0_?q;�0P�K_FI� 	�$THKYGPA�NE�4 � DU/MMY1dDDd!ROE4LA!R�!R��	 � $TI=T�!$I��N ��Dd�Dd �Dc@�D5��F6�F7�F8�F9�G0�G�GJA�E�GbA��E�G1�G �F�G1��G2�BJ1SBN_�CF>"
 8F CNV_J� ; �"�!�_CMNT�$�FLAGS]�C�HEC�8 � EL�LSETUP �� $HO30I�O�0� %�SMA�CRO�RREPR�X� D+�0��R{��T UTOBAC�KU�0 }�)DEVIC�CTI*0�� �0�#��`B�S$INT�ERVALO#IS�P_UNI�O`_�DO>f7uiFR_F�0AIN�1��x�1c�C_WAkd�a�jOFF_O0N.�DEL�hL� ?a8A�a1b?9a�`FC?��P�1E��#�sATB�d�M��MO� �cE �D [M�c��^qR;EV�BILrw!�XI� QrR � � OD�P�q_$NO^PM�"Wp�s�r/"�w@� �u�q�r�0D`S� p E R�D_E�pCq$F�SSBn&$CHK�BD_SE^eAG� G�"$SLOCT_��2=�� V�d¾%��3 a_E�DIm   �S �"��PS�`�(4%$EP�1�1'$OP�0�2�a�p�_OK�UST1P_C� ��d��U �P/LACI4!�Q�x4�( raCOMM� ,0$D����0�`���EOWBn�IGALwLOW� (Kt�"(2�0VARa�Є@�2ao�L�0OUy� ,Kvay��P9S�`�0M_O]��ޗ�CF�t �X� GRP0��M=qNFLI�ܓ�0UIRE��$g"� �SWITCHړA�X_N�PSs"CFu_�G� �� WARNM�`#!�!��qPLI�I�NS]T� COR-0b�FLTRC�TRA�T�PTE�� $A�CC1a�N ��r�$ORI�o"��R�T�P_SFg����CHG�0I���rTא�1�I��T�m���� x� i#�Q��HDERBJ; C,�2'�U3'�4'�5'�6'�U7'�8'�9s!��O`T <F П�����#92��LLEC�y�"MULTI �b�"N��1�!���0�T_}R  4F STY�"�R`�=l�)2`�����`T |� �&$c�Z`d�pb��P�MO�0��TTOӰ�Ew�EXT����ÁB���"�2� ��[0]�}R���b�}� D"}����Q����Q�kc���� �^ȇ1��ÂM���P��� Ƌ� �L�  ���P��`A��$JOBn�/�i��G�TRIG�  d�p�߻���³�7�������J0CO_�M�b! t�pF̝ CNG AiBA � ����M���!���p � �q��0��P[`��,��)�"6���0t�B񉠎"J��_Rz�gC�J��$�?�Jk�D�%C_�;���Б��0h ��R�t#�� ������G|���0NHANC̳'$LGa��B^a��� �D��A�`��gzRɡ�!��p�fDB�RA��AZ�0KELT��Ė��PFCT&�b�F�0�P��SM��cI��1�% ��% ���R��a���� S��&���M 00{�o e#HK~�A^S@������۠�t$�"�6SW�CSXC�)�?!%��p)3��T�$@��PANN�&�AIMG_HE�IGHCr�WIDLI AVT�0��H F_ASPװ��`�EXP�1���CWUST�U��&��
|E\�%�C1NV q_�`�a��' \%1y�`OR�c,"�0gsdk��PO��LBSYI�G��aR%�`좔Psp�m��0k�DBPXW�ORK��(��$OSKP_�`ma��"�<qTRp ) ���P���� �0�3DJ!d/�_CN��R�#� �'PL�S�Q�dD�s�DKA7WAw�'�^A�@NFZpfBD�BU��*�"!PR�S�7�
ЖQ����+� [pr�$1�[$Z���Li9,v?H�3ʠ��-�?�4C��9.�?�4ENEy���� /�?�3J0RE\`��20H��CuRo+$L,C,$i38
�? =KINE@�K!3_D�I�RO�`�� ���ȳqvC��h �F�PAÃ3uR�PRN,�B�MR��U!�u�;CR[@EWM �/SIGN��A� x.q�E�Q-$P���.$Pp 2�/� P7�PT2�PD�u`L���VDBAR@�GO_AW���Jp 8� �DCS�pZ�?CY_ 1���@q1<�Q?fIG2�Z2>fN>�����
�qS�&c}P2 P $���RB?�e�P=hP�wg�QBYl�`gT�+1�THNDG�23���KS�SE|�Q��SBL�Y�cc�TK�rR=L�4 HpZ <���VTOFB�l�FEfA�ǿb�TqSW�5�bDOC���MCS�f�`Z$r�b �H� W0��T�eS�LAV�16�rINP��f��LyqQP�_7� $,�S����=��v��uFI��r줭sc�!���!W1ԭrNTV�'��rV	��uSKIvTE�@W���:�&J_� _�00��SAFE�A�_S}V��EXCLU��*B �PDJ L1�k��Y�d�ƻrI_V<� !PPLY 0b�旁DE~w��_ML�2�B $VRFYi_�#��Mk�IOU@��憻 0���:�O�PƜ�LS�@jb;�35H72��Sr�� Px%�X�{P�hs� �� 8 @� TA� qঠ� 2t_SGN��96����@�A��� ��iPt!��s"��~UN�0jdՔ�U���B �@� ��� ����bl�OGI�2:� @�`Fؒ���O�T�@@�:41(�774�C2�M`NI�2;��R������A�q��D{AY1#LOAD�T�/4~�;30� �EFV�XI�b< @%1�O㠈3� _RT;RQ��= D�`@���Q@  �EjP"�㥎�<�B�� <	�@��AMP��]>�a�����a�8S�q�DU�@q���"C�AB��?A��0NSls���IDI�WRK�h^�� V�WV_]�~��> �DI��q�@� /.�L_SE2�T���/��Z`��0��#�E_п�u�v�j��SW�J�j� 𲰂�	���=�c�OH�z�PPLJ�v�IR!��B� ���w�d��B"����BASh��� X ���V�����?C��Q��R7QDW��MS����AX}�8�u�LIFAE� �7�A1C�NJ� ��S��H���Cs�>�Z�C`QN"䘡U��OV� _�H9E����SUP�hb�C�� _�Ԥ���_P����[Q��Z��W����ו�Tb��XZX$ `1��Y2F�CM@�T��t@�N�p��qpP��9A `�P�.�HE��SIZ�y֥�u��BN�pUFFI���p� �Q�/40�<2671^@�DwMSW9B 8�KEYIMAG�CTM@A��A�Jr||#��OCVIET�N��C C�V L�t<���s?� 	3q� j:D�"pST�!x�0�� 0��Ѡ���0���EMAIL����@����c`_FA�UL��EH�CC�OU�p}$T@��F�< $���eS�]���ITvBUF@��q���T  ���	BdC�t����#��SAVb$)�e� �A� }���Pi�e@U�b`_ H���	#OT{BH�lcPր(0�
{��AX1#��X @��_GJ�
�YN_�� Gj�D��U/0e��M��*��T8�F��ِ�A!H�(@u��&�C_r@�@K�D����=pR���ugDSP �uPC�IMb��J����U��ЁEƀ��IP��su��D`�TH�0�c��TuA�H�SDI�ABSC�ts��0Vzp*} X�$�#��NVW�G�#��$0� FJ�/d0�j�ASC��U·MER��uFBgCMP��tETH��!AI��FU��DU` �a�@;⠂CD��O � ���R_NOwAUTg` J���Pp2��n4ĥPS*m5C`}5CI�.�ak3� =KH *}1Lp��Q� �&�I���4#Q�6s���6ѡ�60��6���67
�98�99�:J��8�:U1J1J1J1+JU18J1EJ1RJ1_J�2mJ2�;J2J2�J2+J28J2EJ2�RJ2_J3mJ3�:3�KJ3J/�G8J3�EJ3RJ3_J4mB�N}�EXT�>aLC`��F�fF�5Q9gܒ5��FDR�MT��VC��C�wa\}"C�REM,�FANj�OVM��eA�ioTROV�iDTm 6�jMX�lIN�i�М�j�IND�`!�
xxp /$DG ���`opS�9�D��`�RIV)0Qbj�GE[AR�IO0�K�bu�Nj�x�.؎��p|�qj�Z_MCM>��C�d`��UR)2N y,{1��? ��r
 ?��H�?�q�E���q0�T0lbO�ߠ��P� �RI�T5��UP2_ gP Ѡ#TD=  ��C����qP�J����C;Q T��$9 ZO�)��OG��%E�8�3e&0IFI��e�0�0����PT���caMR2ieR� vbY�vbLI q��{g����f��Ŗb_mAN~F�_�F�I4+�M;v`r}D�GCLF��DGDMY��LD�q>t5[�P5S�كk�SY�M�? T�FS� l�T P�)���
�/$EX_)�@�)��1�� ��*�3b�5�b��G�!ieU �� p&2SWKO��D�EBUG�S��0�G�RY�zU�#BKUv� O1�@ O�PO8��Π0��Π�MS]�OO��S�M]�Eq؁pQ`_?E V $�X���p�TERM2�W<;����ORIĀ6�yX;�_`�SM_���$7�Y;����TAry�Z;�#��UPB�[� -��Qb�V$G���W$SEyGźאELTO���$USE0NFI����p���`�>��X$UFR����`q0豈�D5h�OT1�ƴ TA_ �C�NSTd�PATT!��Y�OPTHJ!B0En�8�K0�ART� ��p������REL��&SHFTF"�_�.��_SH��M�!B0"x� ��n���Z����OVR
#&SHIԾ���U�2 �AY#LO$ 5I1�p_�d���d�ERV�0 *�} ��b?�d��Q0����A��RC
���ASYMh���WJ�apE�����f�2�U��d�5����D5��P#Gи!	�O5Rd�M���!���\��΢�^��87��k�] �E�]��TOC���q��OP��N z�3�&1���aO�a> R%E��R�#&O0��`�e��R]�����|����e$PWRSp3IM��[�R_����VISy�r���UD��t�� ^>��$H����_ADDR9fH$�Ga�z��s�i1R� =_ H8�S� ��S��C0��C��CSE�a�baHSO0��` $���_D`�v��PR��1wHTT� UTH��a ({0OBJE�1u���$9fLE�P�-=b � �*g!AB_qT���Sk�#DBG�LV5#KRL"�H�IT�BG0LO:���TEM4$�0�b������SS�p�4�JQUERY_FLA��f WYA���ec��� PU�"B�IO0��4G���H��HB �IO�LN~�d/0i�C^��$SL�� oPUT_�$���Pwp�rSLA�� e/2�����ӡ�ҽ1IO F�_AS�f��$L��U���#�04�#0����,�HYOgN!v'$TY!UOP�g ` l!9f�b>$�`E&�!��P����'а!E&�"�&��P_�MEMBk0T 7h X IPz�v��"_#0v����0��pOc6�1w�DSP��' $FOCUSB�Gv��0UJhfi � 60S��JOG��W2DIS�J7z��O��$J8�9�7��I6!�2�77_LABQ����0�8�1oAPHI�pQ�3:�7D+�J7JRA4`�P�_KEYp ��KILMONz�j&`$XR �=0cWATCH_0 �DӘ�U1EL� �1yc`B�k GpG�qVP�-ffBCTR���fB5baLG|�l ���+h�"��LG_SIZ{Y��E
��F,
 �FFD�HI�H�H ��F�HM��F�@���C 5V
�5V
 5V�@5VM�5W�`S)@S����@)Nv1��mx � �� R��4a�PÀU�Qrk�L�S�RDAU�U�EA I���R�PGqH��� BOO~��n� C-"2�I�TGcd��)&REC�-jSCRN)&DeI(#S��RG�� ��cl�!#��b�!	Sa"Wkd!�T!#�JGM�gMNCHL"FN�2�fK�g7PRG�iUF�h	�n�hFWD�hHL/ySTP�jV�hĀ�h,`�hRSgyH!�{&C�Es��!#���g�yUt�g�¬f|@d6#�bG�i4�PO��JzZeEsM�w82�iE]X'TUI�eIP�cw��c���c���` �a����s��Jg��Ka;NO{�ANA"�·�VAI�0zCL�����DCS_HI��������O�����SI)��S'��hI�GN�@��C�aTܮ���DEV�wLLv��a_BU𠪔�oa@�T���$�GEM'9nD�(cѢ��pa@Ѕ�C�!��OS1��2���3��d_����q �T0v-�絡.e�IDX���X-fL�b�STm R�P�Y0���� p$E��C���  ��p��� ��r L*�</��Q(6����6�E�N 6���Jd_ s Y��P$ d�KaD� �MC�R�t �T0CLDP|m ��TRQLI`0��e0x�f�FL>1���_����DUA��LqD������ORGe0 �r���WX�����Y����V�O�u � 	P���uu���Si�Tx���00�ްS�[�RCLMCi����{ɘm[�C0MI��O�v� d�Q6�RQ�0�0�DSTB��Y� 1��{a��AX��@|�� �EXCES�Ҥԑ��M��wA0@�¹�*����x(��_A�ʊ l���t�V�K|�y \*܃2��$MBLI�E��REQUIR�����O��DEB}U_N�ML�M{�zW�.!��B�ӊi���N,03Ѩ�{0�R�RkHV�DCE��T�IN3 `!�TRSMw0p�S�N�����s<��ZA�PST�  �|h�LOC9�RI,� 9�EX��A��:������ODAQo%}���$@�Q΂MF �A�_���p�C���P��SUP�M�F�X��IGG�"~ �0��MQ���v�5@� %����m ���m ����6#DATA����E� 1B1MQ" �N�� t�MD
IF)?�!��H���1!� �1"ANSW�a!ܑS�
!D�)��H3Q�$�� ?�CU�@V0_ >0���LO�P$��=ұ���L2�p�����RR2I5��  ��QA�X� d$CALII��NUG�2g�RINp<$R�SW0��K�A�BC�D_J2SqE����_J3v
p1SP�@6 ��	Pp�3��\�����J���P�O村IM��[�CSKAP��$�P�$J�Q[�Q,6%%6%,'���_AZW��h!ELx�����OCMP�����1X0RT�Q�#�c1�c@�Y�1��(t�0�*Z�$SMG�p�����ERJm�*�IN� ACߒ���5�b��1�_B�542d���14X�͆>9DI~!��DH� �30���$V�o�Y�$�a$�� 
��A���.A ���ňH �$�BELy lH�ACCEL?��8���0�IRC_R��'��ATw�c�$PS �k�LM�yP D���0G�Q�FPAT!H�9WG�3WG3&B��#�_�2�@�AV�
��C;@�0_MG|a�$DD�A@[b$FW(����3�E�3�2��HDE�KPPAB�N.GROTSPE�E�B��_x�,!��D�EFg��1M�$U�SE_��Pz�CD ���YP�0V� �YN��A{`uV�8nuQMOU�ANG�2�@OLGC�TINC ~���B�D���W���ENCS����AX�2��@INk�I&B0e��Z�, VE�P'b23_UI!��9c/LOWL3��pc x��UYfD�p��Y�� ���Uy�C$0 fMOS`���MO����V�PERCH  vcOV�$ �g9��c�� \bYĄ��'�"_Ue@0��A&BuL�������!ec�\jWvrfTRK�%h�AY�sh� �q&B�u�s���&l��Rx�MOM|���h��� ���C�sYC���0DU��BS_BCKLSH_C&B ��P�f�`}S�7��RxB��Q.%CLAL���b?��pX�t�CHKtx�H�S�PRTY��B��e�����_~�N�d_UMl�ĉCуΫASCLބ PLMT�_L�#��H�E������E��H�-��Q#p_��hP	C�a�hH��ЯEǅ�Cw��XT�0�GC�N_(N�þ���S	F�1�iV_RG�e�!p��&B���CATΎSH~�(�D�V���f�'A�	� �@PAL΄�R_Pͅ�s_y��뀎v�`x��s����JaG5�6Ф�G`OG��>�rTORQUQP� �c�y�@�Ңb�q�@�_W�u�t�!�14��3�3��33�I;�II�I�3F�&������@�VC�00��pҩ�1௾2�ÿ�¶�JRK���綒 DBL_�SM�QO�Mm�_D9L�1O�GRV:�3�0�33ģ3�H_��Z@a�COSn˛ n�LN���˲��ĝ0�ɀ� ��e��ʽ̃��Z���f�MY���z��TH��.�THET=0beNK23�3X�l�3��CB]�CB�3C��AS���e����3��]�SB�3��h�'GTS@! QC����'y��'����$DU��;w	��Q������qQ����$NE�$T�I�����)I7${0L�AP�y��`�k�k�LPHn�W�1eW�S���������W���P������{0V��V��T�0��V��V��V��UV��V��V�V�H�����7�����UH��H��H��H�UH�O��O��OF	���O��O��O��O���O��O�O��F�W�}��	�����SPBALANCE��{�LE��H_P�S�P1��1��1��PFULC5\D\���:1��!UTOy_��ĥT1T2��22N���2, ���@�q^<�-B#�qTHp�O~ �1$�INSE9G�2{aREV�{`�aDIFquC91�l('o21�dpOB!d�=��w2��7P���?LCHWARR�2�AB���u$ME�CH��ДQ�!��AX�qPB��&r�~2��� 
�"��1eROB�`CR r�%�����MSK_|�4� P �_OPR�1�2(47Qst1�,`*R(0)cB�(0�|!IN!�MT�COM_C���0��  �@0 �A�$NOREc�2��l ~2� 4�G�R��%FLA!$XYZ_DA��LP;@DEBU�2 X�0lR�0� ($mQwCODS� �2��r� �p$BU�FINDX*P ��2MOR3� H%0�p�0��:@�p�Q8B�"�1��NF��TA9Q"@�2�rG�.B� � $SIMUL���0�As<�AsOBJE3�F�ADJUS�H�@A�Y_I��xD�GO�UTΠ�4�p�P_F-I�Q=8AT#�Y ,`W�1P +�PQ+ t9�uDjPFRI ��PUT0�RO�
`E|+�Sp�OPWO���0�,@SYS�BUi� @$SOP��QBy��ZU�[+ PgRUNn2�UPA;0!D�V�"�Q�`_�@F���PP!AB�!H��@I�MAGS�%0?�Pf!IMQAdIN$���RcRGOVRDEQ�R�@�QP�Pc�� L_��feÂސ�RBߐ<pX�MC�_ED'@�  H�N�i M�bG��MY119F�#@EaSL30�� x $OV�SL�SDIsPD�EXǓ�f֓Hq�bV+��eN�a
��Pp�c�wx�bw��0Ea_�SET�0� @0�Cr�%9�RI�A3��
Vv_��bw{qnqzp#@-!�@� �4ByT� àATUS�$TRCA�@PBN�sBTM�w�qI�Qªd4F��s�`0� �D%0E�P�b�rr�E�1"�qQpd��qEXE�p���a�"��tKs1�Rp&0�pUP�01�s$Q `XNN�w𓱪d���y �PG�|5� $S�UB�q�%xq�q|sJ_MPWAI$�Ps���LO ��1
 �E�$RCVFAIL#_C@1�PÁR%P�0��#���Ȕ� �
�R�_PL|sDBTB8á���PBWD��03UM��IG�Q `�,�TNL ��b�AReQ�2���qP�¤@EǓ��֒��DE�FSP� � L%0� ��_���CƓ�UNI�S�wĐe�RX)��+�_L
 P�q}�qPH_PK�5���2RETRIE�|s�2�R{B���FI~�2� � $��@� 2��0DB�GLV�LOGSCIZ�C� ���U�"2|�D?�g�_T:��!eM�@C
 #EM���R��y0�8CHEC�KS�B�Po01�B�0.�0R!LbNMGKET��@�3砹PV�1� h�`A�Rp� �1)P�2>�S��@OR|sFORM3AT�L�CO�`q�d���$Z��UX�P�!r�LIG�1� w ˣSWIm �6���,�G�AL_ �� $`@��BԈa��CS2D�Q$}E1��J3DƸ�� T�`PDCK��`�!LbCO_J3�����T1׿�3��˰C_Q�` w� ��PAY��,S2u�_1|�2|�ȰJ3�ИˈŬƗ�tQ�TIA4��5��6S2MOMK@������h����y0B׀AD�ð������PU��NR��C���C���?q���4�` I$PIN�u�41�žӁ�:q �R~ȇ��ٯ��:�@h��a�֬��ց�1��'1R\uSPEED G��0�؅��7浔 ؅�%P7�m�F��U��؅SAM =G��87��؅MOV	B� e0�� ��c2��v� �浐�� ���c2nPsR�����İ$QH���IN8�İ��?�[�6�؂�A���X����GAM�M�q�4$GE�T1R@�SDe�mB
��LIBR[�y�I.�7$HI�0_5a@$c2E`@#A@ 1LW^U@	� 1a¬&o�ʱC=�n �S`�p �I_��pPmDòv�ñ'�����mD��	ȳ ��$�� 1�*�0IzpR� DT#|"c���~ LE^141�q�wa�?�|�MSW�FL�MȰSCRk�7�0��Ѻv���Z 0�P�@9@����2�cS_SAV�E_Dkd%]�NOe�C�q^�f� ��u� ��}ɕQ��}���}*m+ ��9��ժ(��D�@�� �������b31�R A�Mam�7
5�#��^����Mtա � F�YL��
A'�VAS	BtRna`7GP�B
B�l3
A%`�GSB1W? �2�2cЬ3oBB1M&@�;CL�8���G$�b�1v���M!LrǢ �N�X0�d$W @�ej@b�� @=� BD�BK�B�-�> @�P����ycİX �	OL�ñZ�E���uԷ� ��OM �R/d/v/�/�/��A��j	�Le�_��� |��H ��jV��yV@��yP�ʗW�V��E�P��8�MS��8����NTP=��PMpQ}U�� � 8Tp�QCOU,�QT�HQ�HOY2`HY�Sa�ES��aUE� `"#�O���  b �P�0�rUN�pʌ3��O$�J0� �P�p^e������O�GRA�qk22�O��d^eITm�aB`INFOI1���k�a�k2��OI�b� =(!SLEQ(��a���`�foaS� ���� 4TpENAB|LBbpPTION|s�����Yw��1sGCF:��O�$J�ñfb���R�x!�]|ot:�OS_EDŀNJ0� �N��@K��j��ES NU�w��xAUT,!�uCO�PY�����v�8 M�N���PRU�T�� �N�pOUN��$Gcbn��a_RGADJI1�2�3X_B0ݒ$ ����@��W��P������@㊀��EX�YCZLB��NS6u�N0άLGO���NY�Q_FREQZ�W`���+�p�\cLAm�"����Ì�uCRE�  c� IF�ѝcNmA��%i�_GmSTATUQPmMAIL�� 1��y�d����!��ELE�M�� �7 DxFEASIGq2��v���q!�er$�  I �`�"��ae�|I��ABUq�E�`D�V֑a�BAS��b� �[�Ub�r % $�y���RMS_TR C�ñj���Ca��ϑ���,r���C�YP	~ � 2� g� �DU�����Ԣ�0-��1��1���qDOUd�ceNrs��PR30z;p�rGRID�a�UsBARS(�TY�Hs��OTO�I1��P`_��!ƀ��l��O�@7t� � �`�@POR�cճ��.ֲSRV��)���DI. T���!���+��+�4)�5)�6J)�7)�8��aF���:q�M`$VAL�U|�%��R��7t�� Cu'!�a��1�� (gpAN#��⛑R�p0� 1TOTcAL��[��PW��It�&�REGEN$�9��SX��sc0��Q����PTR��Z�$�_!S ��9дsV���t���rb�E��x�a�"�^b�p��V_H��DqA�C����S_Y4!��B<�S�AR�@2�� f�IG_S!Ec���˕_b`��#C_����w��?r��8%�b�H�SLG#�I1��p"=���4в�S�2̔DE�U0!Tf.p��TE�@���� !a�����Jv�,"��IL_M`K��z�н@TQ�P��a����2VF�C�T�P���^�Mu�V�1t�V1��2��2���3��3��4��4 ����С���1v�"IN	VIB@PN�; �!B2>2JU3>3J4>4J�I05���"���=p�MC_F`3 � L!!�r��M= I��M� �[PR�� KEEP_HNADD��!f�C�A�� !����"O�Q �I����"��?�"REM9!�ϲ^�uzU��e!HP�WD  S/BMSKG�a	!�B2B�
#COLLAB�!��2����4�o��`IT��A`��D� ,pF�LI@��$SYNT� ;,M�@C>��%пUP_DLYI1�MbDELAm ј�mY�PAD�Ax�`�QSKIPE5� i��``On@NT�1� P_``�b�'�` �B9P�'���)3��)� �)O��*\��*i��*v���*���*9�J2�R‎��?sX��T%�|1�{2ܐ�|1��a��`RDC!F�+ ��pR�sR�PM��'R^��:b�2�R�GE�p2��3d�FL�G�Q�J�t�SPC��c�UM_|0��2/TH2NP�F@o0� 1� �0E�F�p11��� l`[P�E-Ds#ATW o�[�w�B�`�d�A�p3�BfcAHnP�B��
_D2gB�mOO�O�O(�O�O�G3gB��O�O@_ _2_D_��_D4gB�g_y_�_�_�_�_�G5gB��_�_oo,o>o�G6gB�aoso�oP�o�o�o�G7gB��o@�o&8�G8gB�[m����E)S����\@ǡ`C�N�@ �_@wE��^� @o��&m�IO�ፉI���ړ!R�@WE!� W�: �1���0�� �5%Ȃ$DSAB;���֒ �h CL@��­0S232s�̓ ��0�u.��IgCEU{���PEV@>��PARIT�њ��OPB ��FLOW�TR2�҆]����CUN�M�UX�TA���INTEORFAC3�fU����CH�� �t� � ˠE�A$L����OM��A�0"נI���/�A�	TN���Tо ��ߓ��EFA� �"!�Ҏ��� u!��� �O�� &*�� ������  2� ��S�0�`�	�' �$3@}%:B��䎣�_���DSP���JOG��V�h�_P�!s�ONq0%�0����K��_MIR����w�MT7��A�P)�w�>@"���;AS�������;APG7�BRKH����G �µ!! ^���i���P���<����BSOC��w�N���16�SV�GDE_OP%�FSPD_OVR��u �DвӣOR$޷�pN��߶F_���6��OV��SF�<���
�F0����UF�RAF�TOd�LC1Hk"%�OVϴ ��W[ ���8�Ң��͠;�  @ BT�IN����$OFeS��CK��WD����������r���TRr��T�_FD�� �MB_C �B��B����(�.Ѻ�SVe��琄�}#��G)�<�AM��B_0��jթ�_M@�~�x�ቂ��T$CA�����De���HBKX�����IO�������PPA���������Տթ���DVC_DB��?����A���,�X� b��X�3�`���3�0����ϱU8󳠈�CAB�0��ˠ��c� �Ow�U�X��SUBCPU�ˠS�0�0�R�����!�A�R�ł�!$HW_Cg@A��!���F��!�p� � �$�U r�l�e�AT�TRI��y�ˠCY�C����CA���FLT ��������vALP׫CHK�o_SCT��F_e�cF_o����FS�J�j�CHA�1��98I�s�8RSD_!�0���恩�_Tg�7��� �i�EM,��0M"f�T&� @�&�#ޮDIAG��RAOILACN���M�0 �"��1���L���{�PRB�S   ���C4�&�	��F�UNC�"��RI	N�0 "$�7h�� S_��(@��`�0p��`A��CBL� �u�A����D�Ap�a���LD@ܐð�����j���TI%��@�$CE_RIAAV��AF�P=�>#,��D%T2� C��a��;�OIp��DF_aLc�X��@�LML��FA��HRDYO,���RG�HZ 7�����%MULSE�� �����k$J�ۺJ����FAN?_ALMLV�1�WRN5HARD�r��Fk2$SHADOW|��Q��O2 s�0N�r�J�_}����AU- R+�TO_SBR���3���:�e�6�?�3MPIN�F@{��4��3R3EG�N1DG�6C1V��s
�FLW��}m�DAL_NӀ:����B�	����a�vU�$�$Y_B�ґ u�_�z��7� �/�EGe����ð�AAR������2p�G�<�AXE��wROB��RED���WR��c�_�M��S�Y`��Ae�VSWWcRI���FE�STՀP����d��Eg�)�$�D-�{2��BUP��t\V��D��OTO�19)���ARY���R0���6�נFIE����$LINK�!GkTH�R�T_RS���E��QXYZt��Z5�VOFF��b�R�R�X�OB���,8d����9cF�I��Rg��􃻴,��_J$�F�貿S��q0kTu[6��1�w �ad�"�bCԀ+�DU�º�F7�TUR0X#�e�Q�2X$P�ЩgFL�Pd���@p�U�XZ8���� 1�J)�KʠM��F9�p��ӓORQ����fZW30�B�O Pd�,��t����A�t'OVE�q_BM���q ^C�udC�ujB�v�w0L�wg��tAN=�Q �qD!`A�q��=�}��q �u�q���dC��"���SERϡj	�E��HT�ńAs�@�Ue�X��W����AX ��F����N�R�� +��!+�� *�`*��`�*��`*�Rp*�xp*�1 �p*�� '�� 7�� G� � W�� g�� w�� ���� ��� ��đ��DEBU=�$8D3�h����RAB�����r�sV��<� 
�� i�`A��-񷧴���� ��a���a���a��Rq���xqJ$�`D"�R9cL�ABOb�u9�F�G�RO��b=<��B_���AT�I`�0`�����u���1��AND fp�ຄ���U���1ٷ ���0�Q�������PNT$0M�SE�RVE�y@� $�%`dAu�!9�PO��[0ЍP@�o@*��c�x@�  ]$]�TRQ�2
\�d�Bf��j�D"2�{��" � _ � l8"T�c6ERRub��I��VO`Z���TO	QY�V�L�@)�1R��ʄ G;�%�Q�28\�T0e�� ,7��ڙ��]�RA#� O2� d@���[�nq� �Y@$�ph�t � [�OC��f��  ��C�OUNTUQ M�D�SFZN_C;FGe�� 4B�F��Tf4;�~�\� �
��V�}Ѱ�uC� ���M: �"`A��U��q: �FA1 d�?&�X�@=����_B�A<�����AP��o@HE�L@��� }5�`B_BAS�3�RSRF �CSHg�!��1
ש�2��U3��4��5��6���7��8
ל�ROO0�йP�PNLdA�c�ABH�� ��ACK���INn�T��GB$�Uq0� +\�_PUX��@0��OUJ�PH�H���, u��TPFWD_KAR��L@��REGĨ P�P��]QUEJRO �p�`2r>0o1I0������P����6�QSE�M��O��� A�S�TYk�SO: �4D�Iw�E���r!_�TM7CMANRQܨ�PEND�t$�KEYSWITCaH���� HE�`�BEATMW3PE��@LE��]|� U���F>��S�DO/_HOMB O>�_�EF��PR>a9B�ABPx�CO�!��#яOV_M�b[0# I�OCM�d'eQ�}ъ�HKxA� DH�QG��Ue2M�x����cFORCC�WAR�"h�OM>�@ � @r�:#��0UHSP�@1&2�&&3&&4�A��s�O���L"�,�HUN�LO��c4j$ED�t1  �SNP�X_AS��� 0�+@ @��W1$SI=Z�1$VA��տMULTIPL��#! A!� � $��� NS`�B�S�ӂAC���&FRIF�n�S��)R�� NF�ODBU $P���%B3=9G����ny@� x��SI���TE3s�r�cSGL�1T�R$p&�П3a�<P�0STMT1q�3�P�@5VBW�p�4S�HOW�5��SV���_G��� Rp$�PCi�oз��FBZ�PHSP' Av��Eo@VD�0vC�w� ���A00޴ RB% ZG/ ZG9 ZGC �ZG5XI6XI7XI8*XI9XIAXIBXI  ZG3�[F8PZGFXH��TXdI1qI1~I1�IU1�I1�I1�I1�IU1�I1�I1�I1�IU1 Y1Y1Y2WIU2dI2qI2~I2�I2�I�`�X�IQp�X�IU2�I2�I2�I2 Y�2Y2Y�p�hdI3�qI3~I3�I3�I3��I3�I3�I3�I3��I3�I3�I3 Y3�Y3Y4WI4dI4�qI4~I4�I4�I4��I4�I4�I4�I4��I4�I4�I4 Y4�Y4Y5�y5dI5�qI5~I5�I5�I5��I5�I5�I5�I5��I5�I5�I5 Y5�Y5Y6�y6dI6�qI6~I6�I6�I6��I6�I6�I6�I6��I6�I6�I6 Y6�Y6Y7�y7dI7�qI7~I7�I7�I7��I7�I7�I7�I7��I7�I7�I7 Y7jY7Tf�VP� =Uc�� l�נ���
>A820�����RCM2���MbT�R��|���Q_�ЁR-��ń����[�Y�SL�1�� � �%^2��-4�'4��x-Y�BVALU��Ё���)���FJ�ID�_L���HI��I��LE_������$OE�SAb��� h 7�VE_BLCK¡1>'�D_CPU7ɩ  7ɝ �����E����R � � �PW��>�E ��LA��1Saѝî���R?UN_FLG�Ŝ� ����� ���������šH���Ч�}�T�BC2��� � _ B��� br� 8W?�eTDC�����X��3f�S�TH�e�����R>�k�ESERVEX��e®�3�2 �d��� ��X -$��L�ENX��e�Ѕ�RyA��3�LOW_7��d�1��Ҵ2 �MO$/�s%S80t�I��"�`ޱH����]�DEm�41LACE�2�CqCr#"�_MA� pl��|��TCV����|�T�������0B k�)A�|�)AJ��%E�M7���J��B@k�X�|���2p �0:@�q�j�x JK��VK�X�����ы�J0l����JJ��JJ��AAL���������e4��5�Ӵ N1��P ����LF�_�1�� c�CF�"� =`�GROU���1��AN6�C�#\ R�EQUIR��4E�BU�#��8�$Tm�2���|ё �%�� \�APP�R� CA�
$O�PEN�CLOSD<�Sv��	k�
�.�&� �<�MhЫ�8��v"/_MG�9�CD@�C ��DB{RKBNOLDB>�0RTMO_7ӈ$r3J��P��� �����������a6��1�@ � |��%��� �� ���'��-#PATH)'B!8#B!�>#�� � �@�1SCA����8IN��U�CL�]1� C2@UM�(Y"��#�"�����*���*��� PAYL�OA�J2LڠR'_AN`�3L��9�
1�)1CR_F2gLSHi2D4LO4��!H7�#V7�#ACRL_�%�0�'�$��9H���$HC�2�FLEX��J#�� P�4�F߭�����0��� :����|�HG_D����0|���'�F1_A�E �G6�H�Z�l�~���BE����������� �*��X�T,�C���@@�XK�]�o�^Av�T&g�QX>�?��4TX�� �eoX�������������������	-	:J@� �/�M_q�~�۠AT�F�6�E�LHP���s�J� �v� JEoCTR�!��ATN���v|HA_ND_VB��1ܟ�$� $:`F24Cx���SWMs���� $$M ,00�_Y�ni��P\����A��� 3��D��<AM��_AmAA|��NP�_Dm�D|P\ G��E�S�TaM�nM�NDY��� C����0�� >7_A>7Y1�'��d�@i`�P��������"Qs$�� �O�4D'"��J���A'SYMl%A�� l&!��@�-Y1�/_�}8 � �$��� ��/�/�/�/3J	<�:;�1�\:9�D_VI�x�|��V_UNI�����cF1J����䕶� Y<��p5Ǵ�y=6��9 ��?�?>�wc�4�3�a  �$� AS�S  ����s�=�=� h�V�ERSIONp��~��
��I�RTU<�qσ�AA�VM_WRK 2� �� �0  �5�z�������� �	8�)�L�=���!�:�w�^�|�(ܛ݀��7ѭ���������B�SPOS� 1���� < ��A�S�e�w���� ����������+�=� O�a�s����������� ����'9K] o������� �#5GYk} �������/�/1/C/U/ⰑAXgLMT��X#�%�7  dj$INs/�!�i$PRE_EXE��(� �&)0�q��������LARMRE?COV �ɥ"�
�LMDG �����[/LM_IF �ˆ!X/c? u?�?�?�:Q?�?�?�?< OM, 
0�8O��4�cOuO�O�O�NGTOL  ���A   �O�K��{PP)�O ; ?6_,_>_P_{� $BR_�_w�o_�_ �_�_�_�_o�_'oo7o]o�!��O�o�o�o �o�o�o�o+=�Oa�PPLIC�AT��?��� ��J`Han�dlingToo�l �u 
V8.30P/33�@�lt��
88�340�slu
�
F0�q�z=��
2026�tlu���_��7DC3�pJ  ޭsNonelx� �FRA�������B�TI�V�%�s�#��UT/OMOD� E�)�P_CHGAPO�N������ҀOUP�LED 1���� ��"�4�uz_�CUREQ 1���  � >�>��*ސ�4��!��x�=~� ��u���Hm����HTTHKY����w��� 7����%�C�I�[�m� �������ǯٯ3��� �!�?�E�W�i�{��� ����ÿտ/����� ;�A�S�e�wωϛϭ� ����+�����7�=� O�a�s߅ߗߩ߻��� '�����3�9�K�]� o�������#��� ���/�5�G�Y�k�}� ������������ +1CUgy�� ����	'- ?Qcu���� /��/#/)/;/M/ _/q/�/�/�/�/?�/ �/??%?7?I?[?m??��P�TO�@�����DO_CLEAN�܏��CNM  �K >�aOsO�O��O�OD�DSPDR3YRO̅HI��=M@NO_'_9_K_]_o_ �_�_�_�_�_�_�_J�MAX�p�4�1��뇂aX�4"��"���PLUGG���7���WPRC�@B;@?K_�_ebOjb�O��/SEGFӀK�o�g �a;OMO'9K]�o�aLAP�O~Ǔ �������/��A�S�e�w���΃TO�TAL-fVi΃USWENU�`�� ���䏺�P�RGDIS�PMMC�`{qCL�aa@@}r��O�@�f�e��_STR�ING 1	ˋ
_�MĀS���
`�_ITEM1j�  n������ ����Ο�����(� :�L�^�p����������ʯܯI/O �SIGNALd��Tryout �Modek�In�p�Simula�tedo�Out�.�OVERR~�@ = 100n��In cycl�"�o�Prog OAbor8�o���Statusm�	�Heartbea�ti�MH Fa�ul����Aler ���ݿ���%�7�pI�[�m�� �3 f��1x���������� �*�<�N�`�r߄ߖ� �ߺ����������WOR�`f�L���&� t����������� ��(�:�L�^�p���p��������POd� ����d���%7I [m����� ��!3EWi��DEV���� ����//'/9/ K/]/o/�/�/�/�/�/��/�/�/?PALT��81d�?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O&?GRI`f��AP? �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o@o$o6oHo�OR�� �a�OZo�o�o�o�o�o &8J\n��������noPREG<>%��o�L� ^�p���������ʏ܏ � ��$�6�H�Z�l��~�����$ARG�_L�D ?	����ӑ�  	$�W	[�]�����ƐSBN_CONFIG 
ӛ�&�%� �CII�_SAVE  ��E�<�ƐTCE�LLSETUP �Ӛ%  OM�E_IO��%MOV_H�������REP�l���UT_OBACKt�0�FRA:\�� ���_�'`r���=�� J� 	�������ͿĿֿ�6���� 	�1�C�U�g�yϋ�� Ϸ���������ߜ� 5�G�Y�k�}ߏߡ�,� �����������C�U�g�y����a��  )�_�_\A�TBCKCTL.�TMP DATE.D;<��	��-�?�.�INI;0p�8���MESSAG�T�^�_�ېi�ODE�_D��W�8�H���Ox����PAUS���!�ӛ ((O֒��
��*N <r`��������"����TSK  ��=�C�	��UPDT��\�d����XWZD_E�NB\�4��STAp[�ӑ�őXIS&�?UNT 2ӕ`�� � 	S���c2�V0��D�[* Q�����  �`�'$h�
/L/^. "�YK�ާ�J'"��b}��2c/�/_/�/�/�M[ET�`2�P�/�?�/<?�)SCRD�CFG 1C�`��\�\� 1?�?�?�?�?�?�?6��QX��??OQOcOuO �O�O O�O$O�O�O_�_)_;_�O�O���G�R����zS��NA���қ	�wV_[EDZ�1e9�9 ��%-��EDT�-h_ʪ�_o�`/DA���-��_�	�������_�o  ���e2�oɫko�o� 6k�o!hozo�o�c3Y�o��o�n�� 4F�j�c4%�� r���nN��� ����6��c5�a�>����n����̏ޏt���c6 ��-�
�Q��n�Q�����@�Ο�c7����֯ ��n���d�v����c8U��_����0
  }~��0�B�ؿf��c!9!ϑ�nϵ� }J������Ϥ�2φaCR �oį9�K����������n���zP�PNO_�DEL�_xRGE_�UNUSE�_vTI�GALLOW 1��Y~�(*SYSTEM* 3�	$SERV_�GR�R 69���RE�GB�$d� <9�N�UMg��z�PM�U�� 5LAY��  <PMP�AL[��CYC1�0����������ULSU��{�����D��L�N�BOXO{RIk�CUR_;�~z�PMCNV��;�10���T4DLI�4�V���ߨ��'9�K]oR�zPLAL_OUT D�cc�QWD_ABO�R��	��ITR_�RTN���Y� NgONS8� ��CE_RIA_I���<F_1���B =[_P�ARAMGP 1]�w`_�����Cp  �.� � � �� � � � Ȫ � � � �� �  D5`D�$3!g-�<$�H$�T$� DX ʔ X "� B�D1Z� 9X @� 6?� �<HE��ONFI�y���!G_P��1� �e�U? ?0?B?T?f?x?�?�!�KPAUSX�1�UR ,Z��?�? �?�?�?OOOTO>O xObO�O�O�O�O�O�O4_�2O_ey��PCOLLECT�__�Y5auGWE�N��I�"cR QND-EOS�W���1234567890�W�S�u�_��Vy
 H�y) �_#oS��_ohoT�Ao So�owo�o�o�o�o�o �o<+�Oa s������� �\�'�9�K���o��V6Q�2W[ � t>�VIO �YcQyH&�8�J�\��[TR�2؍(�b�
��j��  �x���%�_MOR҂�!� + �'� 	 �5�#�Y�G�}�k����Ӂ"��2A?�!�!3 ҡ�Kڤ*��$R_#*_	�|��C4  AS lyC  x�A3!Oz  BC!�PB/!��PC  @*�����:d�
��IPS$���T���FPROG A%�*6߼�8��I�����&RҴKEY_�TBL  )VR�� �	
��� !"#$%�&'()*+,-�./�W:;<=>�?@ABC��GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~��������������������������������������������������������������������������������͓���������������������������������耇�����������������������1��LCKpۼ3���STA�^д_AUT��O(9��U�INDtTDޞFQR_T1_�Q�T�2��7$����XCƎ 2����P8�
SONY XCg-56�����_�@���u� ���А�HR!5��cT0�B�7T�f�Affrꬿ���� �������5�G�"� k�}�X�����������p��ǼTRL���LETEG��T�_SCREEN ��*kcs�c:U$MMEN�U 1&�)  <���y� �Ã�=& sJ\����� ��'/�/]/4/F/ l/�/|/�/�/�/�/? �/�/ ?Y?0?B?�?f? x?�?�?�?�?O�?�? COO,OyOPObO�O�O �O�O�O�O�O-___ <_u_L_^_�_�_�_�_ �_�_�_)o oo_o6o Ho�olo~o�o�o�o�o �o�oI 2X��hz���� _MA�NUAL�ߕ�DB�L+�DBG_oERRL��'�� �\�n�����NUMLIM�K�d �p�DB�PXWORK 1(�I�ޏ����|&�ŽDBTB_@G )��������qDB_AWA�Y�_�GCP � �=�װ�~�_A!L��D�z��Y��Mt � �_)� 1*�+���
͏�����6�@�_M{�I�SAЉ�@B�P�ON�TIMJ� �ɼp�ƙ
�ۓMO�TNEND߿ڔR�ECORD 10�}� �>�?�G�O����?���2�D� V�h���p������*� ߿�Ϛ���9Ϩ�]� ̿�ϓϥϷ�R���J� ��n�#�5�G�Y���}� �ϡ����������j� ��C��g�y��� ���0���T�	��-� ?���c���\������ ����P�����;�� _q�����(� L%�4[� ����^t� l!/�E/W/i/{// �//�/2/�/�/??��/z�TOLERE�NC��B�В��L����CSS_C�NSTCY 11N6�  ?Β�? �?�?�?�?�?�?OO &O8OJO`OnO�O�O�O�O�O�Oc4DEVI�CE 126� b�*_?_Q_c_u_�_��_�_�_�_�_?�d3HNDGD 36��Cz�^LS 24]�__oqo�o�o�o�o�o�_e2PARAM 5�B��t��dc4SLAVE� 66�e_CF�G 7��gd�MC:\e0L%04d.CSV�ob��c|�r�"A �sCH�p&a&��n��w��f�r��x��ÀJP�>���\_CRC_OU/T 8U����o~EpSGN 9U��Ƣ��\�1�5-OCT-22? 19:30�p��02��4:4�1�p9V UB�u1�݁�nހ��o���Im��P��uG��@uVERSION ���V3.5.1�1E�EFLOGI�C 1:ݫ 	6��|�C���^��PROG_ENBp����͢��ULS{�� ��^�_ACC�LIM|���Xs��WRSTJ�N[���ţ�^�MO�¡Zr,�INIT� ;ݪs5� �*�OPT$p ?	�i�B�
 	Rg575�c��74��56��7��50��R��Ƣ2��6��X�y�TO  ���?�Y�]VP�DEX�d����@W�PATH ;A��A\E������7;IAG_GR�P 2@�k,��"	 E�  �F?h Fx wE?`�D��û ��V1"�ü��T0K��9�Cf�py�pY��dC�pq�B��i�ùmp�4m5 7890?123456��;�����  A��ffA�=qA���pхA��H�Aĩp�������A��Mk����@��tp�p��W0Ae�T0T0�pB4ü� Qô���
���(��A�A�
�=A�L���A���
A�Q�Au��������e������e� Pe�:�د{A�d������dѩp������Au���������r���ߖߨߺ�@�EG��A@�p:�RA5�d�/��)��#P�d�l������"�4�|F�@�Pz�AJ���c�?��9p�A3�\)A,��A&����0���������@�cP�]��AUW�P�J��C���<d�4�-d�%G��(�:�L�^�@��� $HZ��.| ����bt�  2Vh�xm������[���s�����=�
==�G���>�Ĝ��7����8��b�7�7�%�@ʏ�\"&�p�.%��@f�Ah�p9 A���<i��<xn;�=R�=s���=x<�=�~Z��;��%<'��'�~ �?+���C�  <(��U� 4"����&����%ùf��@?Œ?�?@? R?g��$^?�?"?�?�?�?�?�?�?)7L�?S�FB$�/d"Eͽ�>OG��A�Ԭq��sD�L4�x�CA��Gb�tφ���-_7_�C��_����/_�NED  E��  Eh� D�[PbRD_¿�_�86��_�_
z{_�_�w_o�K:o@bù�DP�O=�V��D@66�d��6`���A�U!o�o
o�o��o�o�o�oĿDIC�T_CONFIG; ��Yt؃�eg��ԱSTBF_TTS��
ęVs3���
�iv�[�MAU���Y�M_SW_CF*pB��  �Q�OCVI�EW}pC�}����_�!�3�E�W�i� ;��������ȏڏ� {��"�4�F�X�j��� ������ğ֟����� �0�B�T�f�x���� ����ү������,� >�P�b�t�������� ο��ϓ�(�:�Lϰ^�pς��|RC�sDJ�r!ϐκ��������7�&�[�otSB�L_FAULT �E���xu�GPM�SK_w��pTDI�AG F.y�q��IUD1: �67890123#45��;x�MP�o!� 3�E�W�i�{���� ����������/�A�F�X W!�J�"
�|��vTRECP����
�����M� (:L^p��� ���� $6�]�o�l��UMP_?OPTION_p��F�TR�r`s����PME^u�Y_T�EMP  Èϓ3B�pp �A  �UNI�pau!��vYN_BRK �G�y��EMGDI_STA%�1!�G%NCS#1H�{ ��K��9�/_}d d�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO� �O�O�O�O�I�!�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXo�JO�o�o �o�o�O�o�o+ =Oas���� �����'�9�K� ]�wo���������oۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�o�]��� ����ɏ�����	�� -�?�Q�c�u������� ��Ͽ����)�;� M�g�y��ϕϧ�]�ӯ ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�_�q�{� ������������� �/�A�S�e�w����� ����������+ =Oi�s����� ���'9K ]o������ ��/#/5/G/ak/ }/�/�/��/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OY/KOuO�O�O�/ �/�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oQOcO moo�o�o�O�o�o�o �o!3EWi{ �������� �/��o[oe�w����� �o��я�����+� =�O�a�s��������� ͟ߟ���'�9�S� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�K�9�g�yϋ� ������������	�� -�?�Q�c�u߇ߙ߫� ����������)�C� U�_�q��9�Ϲ��� ������%�7�I�[� m�������������� ��!;�M�Wi{ ������� /ASew�� �����//+/ EO/a/s/�/��/�/ �/�/�/??'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O=/GOYOkO }O�/�O�O�O�O�O�O __1_C_U_g_y_�_ �_�_�_�_�_�_	oo 5O'oQocouo�O�O�o �o�o�o�o); M_q����� ����-o?oI�[� m���o����Ǐُ� ���!�3�E�W�i�{� ������ß՟���� ��7�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���/�9�K� ]�oω��ϥϷ����� �����#�5�G�Y�k� }ߏߡ߳��������� �'��C�U�g��w� �����������	�� -�?�Q�c�u������� ���������1�; M_����� ��%7I[ m������ �)3/E/W/i/� �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?O!/+O =OOOaO{/�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_O#o5oGoYosO eo�o�o�o�o�o�o�o 1CUgy� ������o� -�?�Q�ko}o������ ��Ϗ����)�;� M�_�q���������˟ ݟ�	��%�7�I�[� u��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ�a�� �/�A�S�m�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� e�o��������� �����#�5�G�Y�k� }�������������� ��1C]�Sy� ������	 -?Qcu�������� �$E�NETMODE �1I^��    �(/:+
 RROR�_PROG %�*%}/�)X%TA�BLE  +�h�/�/�/�'X"SE�V_NUM &"?  �!!0�X!_AUTO_ENB  D%#U$w_NO21 J+�9!2  *�*u0�u0�u0�u0(0�+t0�?�?�?N4HI�S3
 G;_AL�M 1K+ �2u< +�?/O@AOSOeOwO�O�?_2.T0  +s1:"��J
 TCP_VE/R !*!u/�O�$EXTLOG_7REQ�6�E9 S�SIZ)_TSTK�FYc5�RTOoL  
Dz�2��A T_BW�D�@�P<6�Q8W_D�I�Q L^�G48$
?"�VSTE�P�_�_
 �POP_�DOh_!FDR_?GRP 1M)B1�d 	�Ofo: W`��������glpw��qŗ��I ����fWc�o�m�o �o�o�o(L7�I�m��zA�P�KA"��>����� 
 E��	�q�@(�C���<�'�`�K�C`}d�C��N��B�y{��F�@UUT��UTF�Ϗj��s���s�OHcEP]���O��#M���*�KA����?��pF��:6:�N�r�9-��z���  �$7@��v�
�������-��+FE�ATURE N�^�P>!H�andlingT�ool � mp�BoEngl�ish Dict�ionary��
PR4D �Stڐard� � ox, A�nalog I/�O�  ct\b�+�gle Shi�ft�  !*�u�to Softw�are Upda�te  fd -�c�matic B�ackup�IF� O��gro�und Edit�ސ�g R6�Camera3�F�7�Part��nr�RndIm���p�shi��ommo�n calib �U���n����Mo�nitor�Ca�lM�tr�Re�liabL��RI�NTData Acquis��Z�ϠC�iagnoqs��0�<�almC��ocument Viewe�\����C�ual Che�ck Safet�y��  - B�E�nhanced �Us��Fr���8� R5�xt. oDIO �fin�s (�@ϲend���Err�Lm� D� p^���s	�E%N�r.�հ �P��rdsFCT�N Menu��v�8���m�FTP ;In'�facN�=��G��p Mask� Exc��gǱi�sp��HT^�Pr�oxy Sv�� � VLOAאig�h-Spe��Sk�iݤ ef.>�H�f�ٰmmunicons�
!�
��urE�'�7�r�t F4�a�c�onnect 2�;�Incr`�st�ru���� Sp�KAREL C�md. L��uaΊ�OAD*�=�Ru�n-TiưEnv�� �D;�(�el u+��s��S/W��.{�Lice'nse����
�����ogBook(S?ystem)蔭��JMACRO�s,��/OffseS�Z�MHٰp���� j73ΰMMRx��l�35.f��echStop��yt�R� ize*�3Mi��O� 2�7��x��0����miz���odM�witc�h����a�.�� yv���Optm���49���filN��ORD��0�g��� 8496�ult�i-T������C�PCM fuyn,��.sv�oO���� �^�5�/Regi��r��	��!2�ri��F� � H59k�1�Nu�m Sel*�  �74 H��İ A�dju���adi�n��O� ,[���t'atub��\У��������RDM R�obot��sco�ve� �d e�m(�ٱn� SW|��Servoٰ�s�ꒄ�SNPX b��1��g P��Libr���1�ڐ 9� ɰW.30g o��tE�ossag� f���@ e����"Lg��/I_�
�I�?TMILIB���~� P Firmn�p��^�F�Acc��x��0���TPTX����510.� el�n���������Hw573�rquM��imula��� �2�Touz�Paxѩ1� T��6����&��ev.��IUSB po�����iP�a�� 0�\sy nexc�ept��3 <� \�h51 ����oduV#��9���Q�VN�k"6PCV�L{&�^}$SP /CSUI�d���+�XC��auҠWeOb Pl���t?  �#S��\"	2��������S�&ު�V?8G�ridplay���&� ��8�-iR�b".� @ � R-�2000iC/1�65¦ d+�+�l�arm Cause/1 ed�<0:ПAscii����L�oad��V4�3Upql�0�_CycL��c�m�ori����F�RA[�am�) t{dt��NRTLi��3Onݐe He�lݨ 542*�P	C`ρ�4�`�]�1�trߵ48��RO_S Ethv�t[�ܿ�10\ҠiR�}$2D PkߵD�ER>1�E����of��A��ΰ�FIm��F��� z��64MB DRAMު�@:��9RFROA[�Ce�ll3� ����shrQ
��Zc���ÍUk�}p� pide�W�tyL�s��|0\$z�!CtdѰ�.��@"oEmai��li����+�\�� R0�q�Z$GigE�N�4OL�@Sup"��b�pW3oa�~�cro�� ����4��QM��Fauest�A>�j�� miH9.dVir�t��W��0{&Im�M�+T���}$Ko�l/ Bui��n�յ'GAPL�&��MyV6�s "�0�*CGP�Yl���{RG�'p�{�SBUW�RQ�)K�&cm\:��z��fXb�)O�võ(TA�&'spoҠ-�B�&���
 I�\E P�+�C�B'fg-��&"�  �E��sv �b��vv�3��S_k���TO;-�EH�f6.:
�E�vfx_z�)�V��tr>�)�hZ%.�F�& � ��r���*�G�&���њr�����H��РJzCTIeAc�pw4�LN�:1�Mr�" #[��Dg�"�M�-�P2��~T�@����vxuIi�-�S�&�S�&��*4�W��2.pc�)VGF��fxw�ʪVP2AU \f1x���N�if�u����"in��VPB^���)��s�D���*�a<s�F�5 �M��s�I��wc�{&Traİ���U,p  ��<���2��RDp	��N��HY���p���-��H���Øp)����� �ϭ����ħ���rдy����í4+�Ϟ�'9L���ӎ��y�9ӫ�yc3�U��B�Oߞq�u��kߍӍ�Sy*�ߩ�\Yyy����k�W�ߞ�ӄ�Yx����:��	�����y��5�o�e/�Q��,�K�m���g��^9~���u�2��A���������F�y�����y�)����|����1�m��.�+�M��8<G�i�7n��c����1�� �����W�����7�{<����6�Z�������uk��[�3|�!��?�ϔ�s�iB\����_F��{�x@.��wrst���B<�� H68���@H)T@J�EE�NDI?��tql[}
_�w�P��TQ (��IG) "���PA�p��T�/��85/A#bs;/�C/U/� ,q�/B�Gp�/�#��/�"36�5�R ?!2Oepai?5!:/pY4W���%INTo? e?_.q�?4)��?�2�pa2g�?�F �O�?A�ad6?��ty ZUD2gunOO�qC533R?�D�0u�O�/�Mcm���OO�LNT�?��P_�����0_QR7�L_�Cfi�._H?_,_f'R50<�_�SAF-F�_�7�w.vo��_�_88�/�dM Cbo����o�bvrEo��p�aa�oaD�@�osF'-AS-sS�p'�Is(�PCesXPL��O�tlo_�ut\�a�Oh%afvh%- B��/����C�$��srp�?@_�?�`w�}�bA�����h��`��]T�ˏ�sg#ch�os�t��CG\s;��us�?���sSg�/�G J��&��GDǟi$"�o�ggdiʏ!�fd��8�?h%J64S��Tut�o�O�?s����F �_����E�0���D`!�)�NO4E�O�fi$II���iwjO�l�ž��>�?*�lb
��V��vjr/��
� ��7��ϥ�_�?zG7\2O�EG��Ϲ?�`��1� ޯ��_d�o�i�8��c�50�>�x�Ͻ�"Lo�h%����dj9�﴿ƿؿ��c� up9�C� #j9{�E��L��Ek,B串����oS_�e_�&/��O}�j94JϬ�duZ��U����=d;�����8���r7�Dhu���;]m T������d��f�a����M����P�-4r 8V��O" #S�d3wc�P�in�`��a�?& HTuR�ef���
�?hcĕg�r"��q.JG	"�erM/��/ ̢/LRA^��uH7�1�/�tCK�/<eT�XP/?i�k1/m5k3.f��riR�ecHG�/�/ cr��NHGRf?L�i�Y�7�hOuX��H\m O��oρ�;H��DD@ �O��*�<�:I�?�?��8d�R�_ hd�g�hgOO�_���gm	h�_h�m��XO�o|O@�O�o�O\/�o0�f�gm�o`��`e۠;iov��yt��"���uR60���#t1mo_�#1��fdr,op7��_����lp>oh���冬~ ߏ�dLgts���&dޏ��/�o�o
�J?<�vr�F���v.R���Ɵpld�56�%4�0�/���reeK�m�X�P)�KCO*O|%56?�OZ� o~����E$io����jߠ���3l ����OR��LcOFvod��_IF��@$�� ߪ�DߦX!B�f Uce��t�4 �&��(M�O�5)e?Ƕ�/���1?Q�D�uk�'�|����`�boto�����-���6�p`�eS ��on*� ��^�lB'����Տ_�8q�_�rdk��4f ��C(ҿȿ¯ԯ�������̟�����
9I��571��t�gadi39Tar��l�ofk�������v3Pa�@� PJ��|*�������f�et�4epg��2�ed�� E�5��RI  �H552� 747��21�pWel/R78�,� ��0ETXJ6�14��ATUP  wmfh G545�p�"6�p�k�VCAM � 7\awC{RI@ ED" G �UIF)!28 { j�CNREM���`�63�a�S�CH  4C �DOCV� CS�Ui�!0 D s�EIOCE�5�4�#R694 w=e!!ESET=S#!�3!�a 73!fanuMASK��?PRXY�_"q7� �0�OCO���"3=P[�#"�ER� J�" 7�!!J�774#!39�  �Eq�G1�LCH� 0#OPLG%J�5000#MHCR�)%PS�17#MCS� 4D"�04 O#J5y5 [#MDSWe!fY1MD#1s#OP#1.#MPR$07�0w"�0�#�  �#PCMX �#R0A�#� & �00�#� ( �&0�$s50( �#PRS� �3J6903FR�D@ 02RMCNny�ndM�93 ~SNBAA��800�@HLB o "Lo�SM�A�0 (Ww"4 on�it#!2  II�)�TC [#TM�ILe �B�`0"K3�@TPA� �Q�TXa�t\j�@E�L�BM250`0/D8���$78�monf�195d SD95\F�UEC 0OP� UFQR@ ��;!C@ \�@�;!O�0pt"VIP��@#� I�@0�!CsSX� �#WEB �#HTT \st2B24 �#CG�Q#{IG�Qtopm�PgPGS!��PRC�@FSH7���w!6( B�8��![�R RBB�- Ci�B01ro�gw!#IF#"09�8-!!` �@�A64:�(AaNVD�!Ld�1h 6a68( c�`�d SR7c!te.p� 0kaч@�bc`� CLI$0?�sb$c9G MS�"5a�` w- A� STY�@wal �@CTO �CJNN0J98�ORS�0G��b��g J�`OL�1A{bn: SENDu�to�!L�Q���@*r�#SLM� 8�"F�VR� MCHN0C9SW!SPBVP�і PL� ds �qV$0�cCCG $p�aKCR�0
Np�QB� �87.f�QK� j�70*`�p�0'3CSnqToo�CTQL���qTB�P�N���@n;pqC�@�Q#�� �p,#�p ��. �%�$07#%� `8D#TmC� QSQ"TE� �[#m� �tTE� g0t"m�P�TTF�Q[�8���@�#CTG�Q�"8���@�#CTH `�T�TI�@#CT'Qe;qs�PCTM�@SC��$0gS��0bod�yqP�@  �<�� �1� 1d��q�aus�a9�H�P[�qW `@06; �GF `8�V@VP2�@ 623R i��@jH?�g� `n�g�B `�" g�D `��g�F�X mna"PVPIH��+ G V�!#V	`o  23�RVK�@,Np�@CV�Q31��934.�vo =R�erne땗�H���i��r���h���A����37� ��"�\srv����b�3b^�- Sr�B"0x���A�J935땼�B�5 (S�O@���g �1�1�R|�j93땷b���EN�5�� aw�m�SK� Lib������� �����	 �"|��h�h�#��b�wm�sk�nE����ql���pyE�  ���!�02�t F�uïբ6ۯm��u�ji-�I&���8 k��8!�Ń�땼P���2�2�2�Mai'�on��_�/r�;pڦh;�;�G��_r؈��!��4\ֶOR�C��+�5�� "T�¦TP��hQ�65�2�1��4���<�xkP�����ߦ�t�P���QrֶSB�� ch_����)�t!0�B�"
̿ h�h땇�;��� c������������x>�Rp� \toֶ�3���cl�W��2 p�"���������� F����b� Qt�a$�϶0t��ܐFsȒ��76�p�t	� A9d���582��ob��|*{�\a��FMQ ���A��migֶ�I�or��wI�j�rfm���Fc���@1�E�YE~� w���R����4�K2Х70r.�E�ld,�lC�� 1PTP]����.�"AD.�F��&3 k���ask���ȍ`4���۳d�ֶے��ER~�7 R�ƫ/�T�?)�e�rv�G?Y?k?}?8�?�?ӹapa��	�d����r�4�M��t�e����79!J�dd/���G�p�ac� T��<6�b�/� QO�&�$vc>�,@Vg��"��eYW��5/�c BJ�h���R5:�d���0�@��I_��raj��e��hQe}�$`��5(Xa�@Ƈ�et榻�1Otd�j��,�_h�\	UI�/k�jo�FO��`�^���F��r��qW6�5q���K �'6ڦu7s W'�b,'��t'?��n��MFR�ֈ;]�lf�ǯ�fr>֛�w�p�/�,@��_U[ǀ�мn�x '_i�{�����O���p`J���[@�o�in7�L�O�9�\^ � R����+mi2״h �j��҇;- f�nt >��MA H�I  H5529ķ (Cߑ21��l?eR78�c��ߒ0AcaJ�614���0A�TUP�����54]5�t-fl�6yE�=�VCAM�tFL?XCRId����o�UIFULX ��28��mo�NREu'��63��WQ���SCH��Cn�DOsCV�gϠCSU1��cxr�0$�;�EIOC%tx\�c��54�oQ��9�T�;�ESET�TeCmo?�S�/��7S��{�MASK��70��PRXY�T�`���7��`�OߐOCO
e�\?�3�ô`>��!0{�?��|�-��oon G?�39!'�ߑõ H82�LCHd��@I�OPLG�tCGM�?�0��GЎ�MHC�R�Go�S�/1_�C�S4�cgm��50�T��?�5$�[���M'DSWMf.�D������OP��X/2L_�PR��K�����{����883n�CM^��0iA,��0����`~�5#�\h88@�+�?�D���.?�*��4��0D�3��o��S4����9��,i�FRDd�/2�E/��MCN5�H�93�K�SNBAv�U"R��HLB�ɃSM�՛ñ�T���Jc52�SaߐTC4��\�TTMIL�e��P���A|�TPyA���TPTX�ŝ5��TEL�ԫ�0䴈P��8�˳���fK�95����95��w888��UECd�wrt �UFRd��__�Cd�2e-�VsCO4��VIP�;��I�TAX~�C�SX�����WEB84����HTT4�kaz��2T�2M/So�yG#��QIG��< .�IPGS=t\rxO�RC��aߐ7�/a��6D�s@>�R7#��!��Oq�� ���P��Ҷ;�A���K�\��$�0 "��4�����NVD4���#�A�dap��8D���68����R7���P��D0��a��o�bܠn. CLI��l\-C���CMS�'���4�d "ްSTY��[�CTOT�tl枱NN����ORSp4�;�1 ��ltiΰOLS�( E���0�T���L��6�@����9@ ��LM4�HV� o�VR���C�S��shc>�PB�V4䫁/�PL�
A�PV��ust>�CcCG4��0nCR�/4 H5��B��z�K�H573����?����\cms��#�st.~TB����! ��7�C�ԓ�?"�awshD?"��I0?"��3��TCd�K�A 4�\sl"EĤpP��� 4�C[П"Ԥ8c��"4�\(��CTF��c���"���CTG�7e3m#G�THd��h� �I��K�CTvC�59m�CTM��5M����Q0��re\g�P���12���04�����%Sv��13MCTWd��9[@_�GFd�SE]�P2d�t+��2�ո� �2d�ell��P%Bd�I���1Dd��a��1F��tap V3PId���CV�!�Vq��UA��CVK��ۣCV#�cor�eL���H"�Hpp!�HK"�Hatc�JH�H�4�I� �IL0H�I�2�H��H+2�IL�Y4=�H���I�e\a�I�2 Z93��I{�H�@NZ+��H �1��K48�Z<A�Ht�{�Il �Z;"�O�Fs \!�Hk"�H{"@o�F[�BPZo�Z���J��Tok �РH��H\��Il�hZ��Z2=[ng-[gToo�I�p�j(��njrobt_�Xbct.�JL� iur�o��I��i�!��F��POz�ling�j��y���Y"r^zۢ�I�p��Geat^j�]��Z��_je�����_��lkҠHm,��H|���Z��A�I  ��_�  ���Gvhm�J{�svnj���H�49\�J�@L�Ij�749{P�Zt\ajNj�@_"g.pj�mcal�0�fu�J��^zhm-��_bg(���o�\ͫ �1�H�! j��;����MT; "�(Cu�zkL��bgft�JlpX����GCT"���Gfyc]�˝26\fߟ�926�l\� Ί�u�>m��;�Mu1l?�Q��7\^�K����7-[˝���_�6�1Nj48.� H�- �H�@R_�L^zi�Pe��K�Я�F8\�}�}�����Ћ� � yRk,�ticMoj+@OoQxs-@�"�3�gCS j+}LB-[�5 HNj+� co�~�L��z��f�k˝lb�jll����-˂��k/�.���LЎ�kwipJ/�on,�Jt\A��8�SK"��� ��uto�o aB������kwm�1 �o��Htp�ʜ �n}��ex-�˝��x����a^jlL�je$�식i��a��/����rej�1��o�Vor�zR����e T�Z[��[GlclN��߭�SOz�̌GZD��to8�{+B�H643N�`�cSG/o��sg�a�Utui��;`�J���`�;�ndm�ndiN�{/�/�/�/�/ �/�/�/??/?A?�?���riΪ! -Kj7950/�n �zk]�895n/�O�t �Z��wsg�K,�>���iag� SG8J�Ю�ogu����KO]Ltw>_@	J6�4�1�s�{F O�>ګcdݛ��`3d_��r-��N74�uy-�3��RINnzlly��(m^���Lܬ��sgc�zI"� #?
+�oߡ\tw/��0.�@�"���(f�_�[y�Kmm�K}�dct^�t]�+�
{PRZWCHK
�k,�;;`y<p��l�K���LN*R852j �@_jR ����tiN�g WJh�ecN�L�F����w�lZ|*�da9t�ʛ�greN���o  S�TD�r7L�ANG�Aoc�e��`��Q�7��R�870�{��8 {(P�ogge�p��!�58\㕏PATTs�� �t9\��c "B�@�V��1�patd���O���������({q㕔�5�a�p[��m�\㕻�7�\aAw��@�a��p6�𫯽�ϯ�gmon���d��0�B�m�@;A��\ ö��K�I��MHCR�51 	H����g\o��@��=R]� H54ۿm�<@E���;!�����Gomm�;a��R�"|�N㕬0F�C��W�P�)Ai6�� Fƫ�\{��itx�#{ ���iaio����D�e6�eve����7C2 R�@RƜPg��7adl��nt��K�RBT�t�OPTN`772'�CTK"'�g�(�x���)� "AZ'�p;q'�q'�tzn&�{ E'�Ama��-� Mu��ncInDPN����<���872��|�d��(��������#���masy��y "M��o��䃲��#et����\p1������\ ��f���lZ ����lp���9���`p��+ V��ail��@?��䇢�䓢��zd�x<�k`��73.f���irdg��- i���e\ ����� S]0j�021"�1W ��(�`�4�� (i6��e,"� "���+���core_�I���l`F��AY��AB��@����H������ABIC��Par;�M�ai�������<� c\�ITX�>���  ����w1��g Jcwlib��Shi�W�4�� t994\�VSSF��� t�t\j9�f "�O�w� t��$%ini�/��pٰ t�p5G�&,� t\vsR&�x�L�%w� tamcylS/+ref.�%$#� tj��%m�� t�[A�&4\z�/�,z�_v�%A�%�a�%_�ol6��l% �%end�/<c?.?@?�R5o[?m>�6�/�dsshf�/+trt�?�<OAE�'F  !`�G��$%��5vi�6<���6 J92�F3���%25 (�%�@e�&�P�%k�4O dn�wzF��T�&`�XEp�n�&g��? nw\�n�?�,nd�V��N�;XnF j���%se�V I/
&�q&Ѹ�U��5r w�%/aF� �F�_�rclR&�0\pw/Y�90�E�o`/"5Of "U<//A+dprm�%g��%�Xrsu/kmS�T_! L`�6/OŔpM�LO��j��nO1|h�ODn�on�|YCwrp�R/�l���E<�Pe\gya��Krgas�o��k��f�v��4x1tf�?m$ra�o�l�a0�omk�_�Tam�N6+�4�`'9K0.Av�Wې�%�@�Ft���XE sV��ДJ7{37�%|*�%�,P��hB "+��Kw�cfF& I����9�98�vtomzFut vV�_	o;�YC����:8\F&�Y/� t0��f��deb^V ��$�0zFؠ"�䠙g���<9\�&��9��Wr}  �su"�s�t�G��X �f� U (�fagn�F PzFlϜ�Via�TX����vd��w��g��HnzF- O�W CH� �$723�F���E(A�ÿտ2蚽Wc�6�WsvF& S�W�J�R6��_�RVo `RV���ӊ��vt��M\etF�XoN�o��Fr��x���+�1T��F?teR� J5�8�O  34	Wg�le,�%,�j�Dq\at"��zFwIta1FlUTA�VϜ�gw��Mad�W�Oa���6d M��e�FT��o90 H�%NT��R69������i;r\ʆMIR��ӊenʆv���F|�3�N�ITCP��Ta0�p���(MM7G�eT^�o \tpʆI��NYBbusJ׈�m� �I�@zFȀ��F������/��W�'g, 0��4`R_(!sw�&s_�YC67\JF��Tf1_����Dfw��W�Ι4achg��a96�_��� _���_r�V�% 9�9YA�e��$�FEAT_ADD ?	������  	 �$YA//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ��߿������DEM�O N�   ��*� �2�_� V�h���������� ����%��.�[�R�d� ���������������� !*WN`�� ������ &SJ\���� ����//"/O/ F/X/�/|/�/�/�/�/ �/�/???K?B?T? �?x?�?�?�?�?�?�? OOOGO>OPO}OtO �O�O�O�O�O�O__ _C_:_L_y_p_�_�_ �_�_�_�_	o oo?o 6oHouolo~o�o�o�o �o�o�o;2D qhz����� ��
�7�.�@�m�d� v�������ƏЏ��� �3�*�<�i�`�r��� ����̟����/� &�8�e�\�n������� ��ȯ�����+�"�4� a�X�j���������Ŀ ����'��0�]�T� fϓϊϜ϶������� ��#��,�Y�P�bߏ� �ߘ߲߼�������� �(�U�L�^���� �����������$� Q�H�Z���~������� ������ MD V�z����� �
I@R v������/ //E/</N/{/r/�/ �/�/�/�/�/??? A?8?J?w?n?�?�?�? �?�?�?O�?O=O4O FOsOjO|O�O�O�O�O �O_�O_9_0_B_o_ f_x_�_�_�_�_�_�_ �_o5o,o>okoboto �o�o�o�o�o�o�o 1(:g^p�� ����� �-�$� 6�c�Z�l��������� Ə����)� �2�_� V�h���������� ���%��.�[�R�d� ~������������� !��*�W�N�`�z��� �������޿��� &�S�J�\�vπϭϤ� ����������"�O� F�X�r�|ߩߠ߲��� �������K�B�T� n�x���������� ���G�>�P�j�t� ������������ C:Lfp�� ����	 ? 6Hbl���� ��/�/;/2/D/ ^/h/�/�/�/�/�/�/ ?�/
?7?.?@?Z?d? �?�?�?�?�?�?�?�? O3O*O<OVO`O�O�O �O�O�O�O�O�O_/_ &_8_R_\_�_�_�_�_ �_�_�_�_�_+o"o4o NoXo�o|o�o�o�o�o �o�o�o'0JT �x������ �#��,�F�P�}�t� ������������� �(�B�L�y�p����� �����ܟ���$� >�H�u�l�~������� �د��� �:�D� q�h�z�������ݿԿ ��
��6�@�m�d� vϣϚϬ�������� ��2�<�i�`�rߟ� �ߨ���������� .�8�e�\�n���� ����������*�4� a�X�j����������� ����&0]T f������� �",YPb� �������/ /(/U/L/^/�/�/�/ �/�/�/�/�/ ??$? Q?H?Z?�?~?�?�?�? �?�?�?�?O OMODO VO�OzO�O�O�O�O�O �O�O__I_@_R__ v_�_�_�_�_�_�_m  h$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲�����������   ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ��������
��	�,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_�oi�$FEAT�_DEMOIN [ d�D`�`},dINDEX9k�Ha�,`ILEC�OMP O�;��zaGb'e�p`SETUP2 �Pze�b��  N �amc_A�P2BCK 1Q~zi  �)hD�o�k%�o`}` Ae�om�o�  ��V�z�!�� E��i�{�
���.�Ï Տd��������*�S� �w������<�џ`� �����+���O�a�� �����8���߯n�� ��'�9�ȯ]�쯁��� "���F�ۿ�|�Ϡ� 5�ĿB�k�����ϳ� ��T���x��߮�C� ��g�y�ߝ�,���P� ���߆���?�Q��� u����:���^��� ���)���M���Z��� ���6�����l��� %7��[���  �D�h��i�`�P�o 2�`*�.VR`� *�c�����JP�C��� FR6�:�.�4/�T X`X/j/�U/�,;`%/<�/�*.FM�/"�	��/<�/<?�+STMG?q?��D]?�=+?�?�+H�?��?�7�?�?�?EO�*GIFOOyO�5eO"O4O�O�*JPG�O�O�5`�O�O�OM_�JSW_Ā_� Sn_+_%
�JavaScri3pt�_�OCS�_o��6�_�_ %Ca�scading �Style Sh�eets0o� 
A�RGNAME.D)T_o��0\so1oГQ�d�o`o�`DISP*�o�o�0�o7��e)q8�o
TPEINS.XMLg�:\{9�aCu�stom Too�lbar��iPA?SSWORD.�?FRS:\��� %Passw�ord Config@��������� ��r�����=�̏ a�s����&���J�\� 񟀟����K�ڟo� ������4�ɯX���� ��#���G�֯�}�� ��0���׿f������ 1���U��yϋ�ϯ� >���b�t�	ߘ�-߼� &�c��χ�߽߫�L� ��p����;���_� �� ��$��H���� ~����7�I���m��� ����2���V���z��� !��E��>{
� .��d��/ �S�w�< �`�/�+/�O/ a/��//�/�/J/�/ n/?�/�/9?�/]?�/ V?�?"?�?F?�?�?|? O�?5OGO�?kO�?�O O0O�OTO�OxO�O_ �OC_�Og_y__�_,_ �_�_b_�_�_o�_�_ Qo�_uoono�o:o�o ^o�o�o)�oM_ �o��6H�l ���7��[��� �� ���D�ُ�z�� ��3�ԏi������ ��ßR��v����� A�Пe�w����*����N�`���֦�$FI�LE_DGBCK� 1Q������ (� �)
SUMM?ARY.DG����OMD:3�s����Diag Su�mmaryt���
CONSLOGi��L�^�������Co�nsole lo�g����	TPACCN�R�%:�wς��TP Acco�untinρ��FR6:IPKD?MP.ZIP�ϯ��
���σ���Exc?eption ߱��_�MEMCHEC�Km�Կb����M�emory Da�ta��֦LN�=)n�RIPE�\߸n���%�� �Packet L�Ϻ��$SA���S�TAT�����ߋ�� %�Sta�tus��<�	FTAP����r������mment TB�D��� =�)ETHERNEU����B�S�����Et�hern(��fi�gura߇���DCSVRF���������� verify all�٣M(��DIFF����/diff�PB���CHGD1�x�� �FQ&���	2��� 5�YGD3p���'/ ��N/�UPDAT�ES.m S/��FORS:\k/�-���Updates �List�/��PS�RBWLD.CM��/���"�/�/�P�S_ROBOWEyL1���:GIG����?/�?��Gig�E ��nosti�c*�ܢN�>�)}�1HADOW�?��?�?5O��Sha�dow Chan�ge��٤&8+�2NOTI��O"O��O��Notif�ic��\O٥O�A��_��2_կ?_h_ ���__�_�_Q_�_u_ 
oo�_@o�_dovoo �o)o�oMo�o�o�o �o<N�or�� 7�[���&�� J��W������3�ȏ ڏi�����"�4�ÏX� �|������A�֟e� ����0���T�f��� �������O��s�� ���>�ͯb��o��� '���K��򿁿ϥ� :�L�ۿp����Ϧ�5� ��Y���}���$߳�H� ��l�~�ߢ�1����� g��ߋ� �2���V��� z�	���?���c��� 
���.���R�d�����������$FIL�E_� PR� �����������MDONL�Y 1Q����� 
 �)�@_�VDAEXTP.�ZZZ��p�G�L�6%NO Ba�ck file <!��U3�M�� 7����G�&� J\����E �i�/�4/�X/ �e/�//�/A/�/�/ w/?�/0?B?�/f?�/ �?�?+?�?O?�?s?�? O�?>O�?bOtOO�O 'O�O�O]O�O�O_(_~��VISBCK��|��*.VD)_|s_�@FR:\BP�ION\DATA�\^_R�@Vision VDt �_�O�_�__o_Ao �_Rowoo�o*o�o�o `o�o�o�o�oO�o s�@�8�\� ��'��K�]���� ���4�F�ۏj���� ̏5�ďY��j���� ��B�ן�x����1����ҟg���MR2_�GRP 1R����C4  B�O�	 
������/E�� ֯�r����OHcEP]���O��#M��^
�KA���?��&�r���:6:�N�R�9-�<Z��A�  v����BH��C`}dC���N��B�{���r���пὫ�@UUT��U�����/Ϫ�>��>c���>rа=����>i�=����>����:���:��:�/:6)�:��~ϗ�2ϔ��ϸ�������z�_CFG� S��T � �a�s߅�0[NO {��
F0��� ��/\RM_CHKTYP  ���O����������O=M��_MIN��L�g�����X���SSB7�T�� ��5�L�,�U��g���TP_DEF'_OW��L�����IRCOM�Ѝ���$GENOVRD�_DO��	��T[HR�� d��d��o_ENB�� ��/RAVC��U�UQ �Υm�X��|��������� �� �OU��[���O����⾥8��:���
,.  C�x �h�������B�ϡ������n�!�SMT'�\�.���+�w�$HO�STC7�1]K[��Y��� MC�L��MI��  27.0�1�  e}�� � /*�1/C/U/g/��!/#	anonymous�/�/�/��/�/? L��8 ;{}/j?��?�?�? �?�?/�?OO0OS? �?�/xO�O�O�O�O? UO+?=?_QOs?1_b_ t_�_�_�?�_�_�_�_ o'_]OoOLo^opo�o �o�O�O�O_o G_ $6HZl�_�� ����o1o� �2� D�V�h��o�o�o��� ԏ��
��.�uR� d�v�������?��� ����*�q������� ����ݏ��̯ޯ�� I�&�8�J�\�n���ǟ ٟ��ȿڿ���E�W� i�F�}�jϱ��Ϡϲ� �ϋ�������0�S� Tߛ�xߊߜ߮���� �+�=�?��s�P�b� t����ϼ������� �'�]�o�L�^�p������/ENT 1=^�� P!���  ������ *��Nr5~Y ������8 �\1�U�y �����4/�X/ /|/?/�/c/�/�/�/ �/�/?�/B??N?)? w?�?_?�?�?�?�?O �?,O�?ObO%O�OIO��OmJQUICCA0�O�O�O_�D1_�O�OV_�D2W_3_E_��_!ROUTE�R�_�_�_�_!P�CJOG�_�_!�192.168�.0.10�O�CC�AMPRTGo#o!�7e1@`noUfRT��_ro�o�o��NAM�E !��!R�OBO`o�oS_C�FG 1]�� ��Aut�o-starte�d��FTP�� ~q���F���� ����9�K�]�o�� ��&���ɏۏ����� Wi{X����o��� ��ğ֟������0� B�e��x��������� ү�������Q�>��� b�t�������q�ο� ���9���L�^�p� �ϔϦ�������%� �Y�6�H�Z�l�3ϐ� �ߴ�������}��� � 2�D�V�h�������� �������
��.�@� �d�v���������Q� ����*<��� ���������� ���8J\n� �%�����E Wi{}O/��/�/ �/�/�/��/??0? B?e/�/x?�?�?�?�? �?/+/=/�?Q?>O�/ bOtO�O�O�Oq?�O�O �O_'O(_�OL_^_p_��_�_(�`_ERR� _z�_�VPDUSIZ  9P�^S@��T>�UW�RD ?EuA��  guest3V$o6oHoZo�lo~o�dSCD_GROUP 3`E|� Iq?YM ��nCON�nTAS��nL��nAXP�n_�E�o9P�n�RTT�P_AUTH 1�a�[ <!i?Pendan�g�~�@}9PJ�!KAREL:*���}�KC����p�VISION SCET�`E��I�!\� J�t��s�����������Ώ��-���dtCT_RL b�]~��9Q
@<FF�F9E39�DF�RS:DEFAU�LT��FAN�UC Web Server����bv odL��'�9�K�]��o��TWR_�`FI�G c�e��R���QIDL_�CPU_PC�9QB�@� BH�ǥMINҬ�a�GNR_IO�Q�R9P��XɠNPT_SI�M_DO�!�S�TAL_SCRN�� �y�+�TPM?ODNTOLY�!���RTY8��&�9�.hpENBY��cƣOLNK 1d�[�`�����1�C�|U�ͲMASTE����&�OSLAV�E e�_˴jqO�_CFGsϦ�UO�D��Ϩ�CYCLE��Ϧļ�_ASG s1f���Q
 W� 9�K�]�o߁ߓߥ߷� ���������#�_��GNUM�S�b�U
���IPCH��j�O_RTRY_CN���Z��U�_UPD�S���U �����g�θ`��`ɠP�_MEMBERSg 2h��` $�e��>��HyɠS�DT_ISOLC�  ���r�\J_23_DS��q�~��OBPROC��n%�JOG�d1i���89Pd8G�?�.���.�?�?�?OQNs��V ����3W~�����������POS�RE��$�KANJ�I_m�K�i�pMON j�k~�9Ry����//�^$�r��k����9%Th��p_L�I�l�k�EYLOGGINʴ��`����U��$LANGUAGgE �����Y �!�QLG��lq��9R��9Px�p� � ��砬9P'�03X�k���M�C:\RSCH\�00\��� N_D?ISP m��DpAMK�SLOCw��آDz ��A�#O�GBOOK n���9P~��1�1�0X�9O%O7OIO[O�mN�Mɱ���I��	��5Ib�5�O�O�5��2_BUFF 1-oؽ�O2A5!_ �2��=_?7Y_k_�_�_ �_�_�_�_o�_o:o 1oCoUogo�o�o�o�o�e4��DCS q>�= =��͏L�O�-�1CUg���bI�O 1r� ��s20���� ����1�A�S�e� y���������я���@	��+�=�Q�|uE�TMl�d����Ο �����(�:�L�^� p���������ʯܯ�p ���7�SEV��u={�TYPl����z�����!�PRS����/S��FL 1s�}����$��6�H�Z�l�~ϯ�TP� l�i��=NGN�AM��A5�"e4UP�Sm0GI��\!�����_LOAD��G� %u:%PL�ACi�2�3�MAXUALRMI�c�W�T���_PR���h�3�R�Cp0t�9��M���3Eݗ���P �2u�� �1V	Zi�00���� ��1��.�g�xU� ����������� ��8�J�-�n�Y���u� ����������" F1jM_��� ����	B% 7xc����� ��/�/P/;/t/ _/�/�/�/�/�/�/�/ �/(??L?7?p?�?e? �?�?�?�?�? O�?$O OHOZO=O~OiO�OK��D_LDXDIS�A����zsMEMO�_AP��E ?��
 b��I�O _"_4_F_X_j_|_RпISC 1v�� ��O�_ ���_�_��Ooo@o�_C_M?STR w:�_e�SCD 1x�M� 4o�o0o�o�o�o�o P;t_�� �������:� %�^�I���m������ ܏Ǐ ��$��4�Z� E�~�i�����Ɵ��� ՟� ��D�/�h�S� ��w���¯���ѯ
� ��.��R�=�O���s� ����п����߿�*� �N�9�r�]ϖρϺ��PoMKCFG �ynm����LTAR�M_��z������и���6�>�s�MEgTPU�ӫІ�vi�ND��ADCOLxXի�c�CMNTy�s l�g` {nn���-�&�����l�PO�SCF����PR�PM����STw�1�|�[ 4@�P<#�
g��g�w�� c���������� ���G�)�;�}�_�q������������l�SI�NG_CHK  �|�$MODAQ��}�σW��#DE�V 	�Z	M�C:WHSIZE��M�P�#TASK� %�Z%$12�3456789 ���!TRIG +1~�]l�U%�\!��S
K.�S�YP�69"EM_�INF 1�� `)�AT&FV0E0�X�)�E0V�1&A3&B1&�D2&S0&C1�S0=�)ATZ�#/
$H'/O/�Cw/(A/�/b/�/�/�/? �&?�� �/�?3/�?�/�?�? �/�?�?"O4OOXO? ?�OA?S?e?�O�?�? _CO0_�O�?f_!_�_ q_�_�_sO�_�O�O�O �O>o�Obo�_so�oK_ �owo�o�o�o�_�_ L�_o#o��Yo� ���o$��H�/� l�~�1��Ugy� ��� �2�i�V�	�z��5�������ԟPNIwTOR��G ?k�   	EX�EC1���2�3��4�5�� �7*�8�9����� �����(���4���@� ��L���X���d���p����|���2��2��2���2��2��2Ũ2�Ѩ2ݨ2�2��3ʉ�3��3(�#R_�GRP_SV 1݀� (�ſ1�x�>Ka����?|�ӣR��_Ds����PL_NAME !����!Def�ault Per�sonality� (from FwD) ��RR2��� 1�L6(L�?����	l d��nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲�����B2]���*�<�N�`� r����<���� ������,�>�P�b��t�����BJ � �\  ��  �����  A�  B��UT��� 
����~���  �������B��p��� � CH CH P �Ez  E�� E�` E��;%�Z��*� �  E���F�@&�U�T Ai�  dx�H�x�	$�Hxd�dڭ� }`(d��8�(xx$$ y Xtd D (DDdpWwX� �	X�vXHX����/y�y (�� !��  7%E	��Em�Xw�$%XH$%P��  �/�/�/�/�/�/??�+?=?O?a?s=F��r?�?�?�?�6��E�2ExB�2
�������?Kزd��'O9NO\OjG��0��|M��ն'4� � W%8�O�O�N �0�G��O�JA  A��C�����_�OC_9W�
  � TB�LY��
��_�\��Q�Y=�C�و�V�`HR0� ʒ_P( @7%?���a�Q?ذaر@��6�&س��2n;��	lb	  ����p�X��U�M`��X � � ��, �rb��K��l,K���K���2KI+�KG�0�K �U�L�2o�E	O�n��@6�@ t�@�X@I��b`�o��C�N����
���}v��#���` q�m�|�kQ?�
=ô��  �Hq�o`!b���9�  ���a� �� ���ذa�s�G��}2�m��o�q��v�O���E	'� �� 0�I� ��  � Q�J:��ÈT�È=��9�l���@|��� }~�Q����R������N8���  '���ap?��P�b!p�b){�B���?�CIpB  X���ذ��C�A�g	���o�P�IB P��8�@����P��ԕرD  �O���O��A�,����Š
�`l�1�?	 ٠p���� p` l`:GT � �t�?�ff0{O��įV� �P��`���a�!�/�?Y)RI�a4�(ذ]�Pf�����a\c\dƃ?33�3-d���;�x5�;��0;�i�;�du;�t�<!�+}�oݯ��b��Sb�P?fff�?��?&�9�@׿�A#$�@�o[,ž�x�	�&f 6�ed�g���Hd� �ϣ����� ���$���H�Z�E�~߾�&eF ��mߺ�i���U���y�X��2���E�0�� ��y�d������� ������?�*�܏r� 8�.o�ߺ����T� );ڿPb���������P��A1��T C�=0�ϵ��Y}��2��������C��W��C�= �` Ca�������(!��`�<���bC@�_;C9�B�A�Q�>�V{È�����Y�uü���
/���Q���hQ�A��B=�
?h����/iP��W���ÈK�B/
�=����Ɗ�=�K�=�J6�XK�r#H��Y
H}��A��1�L�jL�K���H:��HK��/�0	bL �2�J��8H���H+UZBu �a?�/^?�?�?�?�? �?�?O�?O9O$O]O HO�OlO�O�O�O�O�O �O�O#__G_2_k_V_ {_�_�_�_�_�_�_o �_1oo.ogoRo�ovo �o�o�o�o�o	�o- Q<u`��� ������;�&��K�q�\�����Gϭ<���� C�aɏ� Ĉ����C'VF�����+b�����Kc�f�� 
E����T�ٟ�=(��_�h۟��������N��x�����3lC�(��:�H���T�f��t�.3��}�����k���q'�3�JJ�����گ����4�"�]P̲Pf�������⟛�ſ���Ի����/���?�{?�N�u�  fUh�*ϳϞ����π�Ϣ�t�.��R�@���X�bߘ߆ߨ�)Z��ߺ�  ( 5�	������B�0��f�t�  2 E�%p"E[@��NŰ"BC��%@ߏ��%�������)�;��� ����������%n�n�%��%��9Xc
 ��! 3EWi{��������b*[���P�I�v�$�MSKCFMAP�  ��� ^�����pD�ONREL  �X�[��DEX_CFENB�
Y��FNC��JOGOVLIM��d��dDKEY��%_PA�N�""DRUN��+SFSPD�TYw����SI�GN��T1MO�T��D_CE_GRP 1���[\���/��? &?��?Q??u?,?j? �?b?�?�?�?O�?)O ;O�?_OO�O�OLO�O pO�O�O�O_%__I_� _m__f_�_O�DQ?Z_EDIT�$U�TCOM_CF/G 1�Q�_�o"o
�Q_ARC�_�X��T_M�N_MOD���$��UAP_CP�LFo�NOCHE�CK ?Q W����o�o�o�o '9K]o������vNO_?WAIT_L�'�W6� NT�Q�Q����_ERR�!29�Q��� �_t�������*��Ώ�d�``OI��P�x  ��W�_���8�?��4�����B�_PARAMJ��Q���	�����s��� =��345678901��� � ��?�Q�-�]�����u�0��ϯ����������7�ODRDS�PEc�&�OFFS?ET_CAR�PKo�m�DISz�K�PE?N_FILE���!�$a�V<`OPTIO�N_IO
/!аM_PRG %Q�%$*	�ά�WO_RK ��'�� ��K�7U��h��f�(�f�	 a���f�7���M��RG_DSBL  Q�����L�RIENTTO* ��C���Z��M��UT_SIM_D�طX+M�VQ�LCT �%��R_�x$aQ�'�_PEXh`ܜ�b�RAThg d�b�r�UP )�5� � �����X������$��2�#��L6(L?}��	l d'� O�a�s������� ������'�9�K�]�@o���������H�2>� ����/ASew�N�<����� ��1CUg�yH���P��� �  �� � �U�A�  B���PB�����H��  ����U�B�p�������N�P E�z  E�� E_�` E��;(�����Z�/�~��  E��''l���@#���T�AJ(��E!Y! a!)!m!Y!u)%)!Y!(E!�%E!ڎ$�^$A! �	!E!a!�%%	-Y! Y%�-58�Z 99HU%E!�D!	$D%% E!Q481X291�%�)95 �/W#95)%91m5a!�5)/Z7��Z (�8�1a�<a1 EE	�(�Em�494X6E9=8)%E15�� |O�O �O�O�O�O�O�O__80_B_T]F�S_y_ �_�_�Vh�����_�[��%�on�_=o�Kg�]�]&�'4 � W%po�oX� g��g�o�j�A�A��c������o�o$w���tB�(~�`��r�|B�� q�y�$�O���1�'k�'ۆ�3�`��0���P�( @ED�D��q?�Q�C�Z7}��o  �;�	lD�	u� ����p�X�[�2���X � � ��, �W��`H���9H�H���H`�H^?yH�R�l����_�����`C#�B�� C4ӄ����c��9���
=���� �������cBz��Β=a�m�另b �s�� �q���g䟒�챏Ǒ�ٖ�o����e	'� � ��I� � � �q<�=��q�9�K���@a�@g�b����������Ƞ����N��  !'۰��Ɓ"�B�Ղ���т6��� � � ��C�a��	m�~��p=�Bp���@�����px����D� �o޿�o��&��o��5�Ю`Q��?	 ٠U�f� U� Q�:���#�}���?�ff\o�ϩ�;� �p����b"�8� ��?Y
rI��q=�(� B�PK��fɆ�A�A���?33�3��m�;�x5�;��0;�i�;�du;�t�<!��y������t����r�p?fff�?x�?&���@׿�A#	�@�o[�	]���� ��uI��wh���-��� ����������	��� -�?�*�c�u�L��������4�V�X����EjPf��^I� m���� � $��W���� ���9��/ /�� 5/G/�z/e/�/�/�/�/�`�A��$�t�/ C�/"?�(d��>�?��Pn?�/�?}?���(��W�?C�@�` CT��?��j4�j0i1A@I��!���bC@_�;C9�B�A�Q�>V�`.È����Y��uü���
�?�3��Q���hQ�A�B=�
?h��iO�Jp��W���ÈK�B/
=�����Ɗ=��=K�=�J6�XK�r#H�Y�
H}��A��1�=L�jL�K���H:?��HK��O�@�	bL �2J���8H��H+UZBu�? F_�OC_|_g_�_�_�_ �_�_�_�_o	oBo-o foQo�ouo�o�o�o�o �o�o,P;` �q������ ���L�7�p�[��� �����ȏ�ُ��� 6�!�Z�E�~�i�{��� ��؟ß��� ��0�pV�A�z�e�Gϭ����� C�a�/�� �Ĉ��ЯׯCVF�����üKG�j����KH�K�� �
Ep�s�9���90(�91�_�h��y��y��i��N���<�T�3lC����-¢�9�Kϰt?�.3��}e�w��k���q'�3�JJ�͑��Ͽ���P����B5P��PK�Zgt�ǿ�ߪߕ��߹����������$�{$�3�Z�  fUM�����������Y��7�%��`=�G�}�k���)Z�����  ( 5� � ������'K�Y  2 E%�pIFE[@tN�bIFB�!�!� C��0	� T�@į��� �*H3��T fx��T�T�E94��T�D=4H;
 �//*/ </N/`/r/�/�/�/�/`�/�/�/GJ@2��5��I�v�$PA�RAM_MENU� ?����  D�EFPULS���	WAITTMO{UTT;RCVg?� SHELL�_WRK.$CU�R_STYL����<OPT��?P�TB�?�2C�?R_DECSN_0<�L 	OO-OVOQOcOuO�O �O�O�O�O�O�O_._�)1SSREL_IOD  ��Y�=U�USE_PROG %8:%*_�_>SCCRk0ORY@3�W�_HOST !F8:!�T�_�ZT\��_ c�_�Qc<o�[_TIMEi2OV�U�)0GDEBUG�MP8;>SGINP_�FLMS`�gn�hT�R�o�gPGA�` 2�lC�kCH�o�h�TYPE5<A )_#_Y�}��� ������1�Z� U�g�y���������� ���	�2�-�?�Q�z� u�������ϟ�
���eWORD ?	�8;
 	PR<�`U�MAI@��gSU�1E�TE#`�U��	�4R�CO�LS�n���vTRA�CECTL 1�v��B1 I�7 8�W d�ެ���DT Q�����РD � *�����W.��.��P.��`.��"��U	�
���2�:�B�B��*�"���;�S�3�:�B�J��+�=�O�a�s� ��������Ϳ߾��K� a��[ÑĠϲ���� �9�������	��-� ?�̨ߺ�����P�b� L�~ߐؓ���)�;� �'�Y�k�}�oρϛ� �����������+� =�O�a�s��������� ������'9K ]o�0\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz�uX�� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲��ߚ�� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p���� ��� $6H Zl~����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OA��$PGTRACELEN  A�  ���@�$F_UP �����SA�[@?AT@$A_C�FG �SET=CAT@��D�D��O�G6@�OhBDEF�SPD �sL�A6@�$@H_C�ONFIG �\SE;C @@5dT�3B AQaP�D�A1Q@�$@�INk@TRL əsM�A8�EFQPEv�E�W�SA��DQ�ILIDlC��sM	�TGRP 1՟Yb@lAC%�  ��l�AA��;H�N��R�A!PD	� a3C	\T�Ai�)iQP� 	 ��O4VGgCo ´|c^oGkB`�a�opo��o�o�o�o�b"�Bz�o7I~3� <}�<�oN�J���� �f�)��9�_�J�"`z����@
t��� d�ŏ�֏���3�� W�B�{�f�x�����՟������J)@)
�V7.10bet�a1�F @��@�A&�ff�Q2�CPC��`�D�Dk`[�C��T��@ DĠ� Dr� �QBH��`�L��PC5R �A?�  ��CCx����b��P!P��A,����Ap�B�b!P�A1������
�?L��?333Aq@��"��Fff.���b�w:�7��AeC�QKNOW_M  �E{F�T�SV �Z (R�C������ʿ��@ٿ�$�A!m�SM�S]�[ �B�	�E?���Ϗ�T̓E`��2�E@��2�������� L�MUR�S�Y�T�j���AC5����e@�Rۚ]{ST�Q1 1�SKO
 4�U��A�� �߰E��*��߽���� ���J�)�;�M�_�q� ������������@F�%�7�|��Ep�2{�9��A�<������P3��������p�4 ��+p�5HZl~p�6�����p�7� $p�8�ASewp�MAD�0F [Fp�OVL/D  SK�ϼO�r�PARNUM � /�O//T_S+CH� [E
}'F!8�)=C�%UPDF/X)��/3Tp�_CMP_0O�0@T@@'{E�$�ER_CHK50yH!6
?;RS�]���Q_MO�o?�5_�k?��_RES_GzФ~ݍ��?�OO�? %OO*O[ONOOrO�O �O�O�O�O�O��3���<�?_�5��(_G_ L_�3G g_�_�_�3�  �_�_�_�3� �_o	o �3@$oCoHo�3�cox�o�o�2V 1�~�|�1e�@c?��2THR_INR�0�!7³5d�fMASmS ZwMN�5sMON_QUEUE �~�f��0V�� �4N0UH1qNEv6;�pEND�q�?�yEXE��u� �BE�p��sOPT�IO�w�;�pPROGRAM %hz�%�p�ol/�rTA�SK_I��~OCFG �h/\�^��DATARè��@��2����� #�5�G��k�}��������^�ן������IWNFORé܍�wt ȟe�w���������ѯ �����+�=�O�a� s���������Ϳ(�4���܌ �I��� K�_�����T��ENB� ͻ1>ƽ�I���G��2�� �P(O�ҡϳ� ������_EDIT �����>��WERFL�x�c�m�RGADJ M�8�AС�i�?�0�t�
qLֈq���5?�?�!��'<@��*�%���0@�#ߊ��2���F�+	Hpl�G�b���>��A�d�t]$I�*X�/Z� **:c�0V�h�@���Ǟ���B����� ������������ ��b���L�B�T��� x���������:���� $,�Pb�� �����~ (:h^p��� ���V/ //@/6/ H/�/l/~/�/�/�/.? �/�/?? ?�?D?V? �?z?�?O�?�?�?�? �?rOO.O\OROdO�O �O�O�O�O�OJ_�O_ 4_*_<_�_`_r_�_�_ �_"o�_�_ooo�f	���o�p�o�o�dJ� �oL��o#�oGY��PREF �����p�p
L�IOR�ITY����P�M�PDSP�>ߴwU�Tz�4�K�ODUC-Tw�8�\�;OG�_TG;�|�����rTOENT �1��� (!?AF_INE�pp�~{�!tcp{�>��!ud��ˎ?!icm������rXY�Ӵ����q)� p�/�A��p�)�j�M�Y���}� �������ן���8�@J�1�n�U�����*�s��Ӷ}}�����,�>W�%�jfp�/z�H֯K�,������A��?,  �p��������ʿ�u"�ut��}�sF�P�PORT�_NUM�s�p��P�_CART�REP�p��|�SK�STA�w K�L�GSm���������pUnothingϿ������c{�t�TEMP �����ke��_a_?seiban0C� ,S�y�dߝ߈��߬� ����	����?�*�c� N��r�������� ���)��M�8�q�\� n������������� ��#I4mX�| ������3>��VERSI�p ��d dis�abled>SA�VE ��	�2600H721:&�!;���̏� 	(�rmoN+	E/`�eb/�/�/�/D�/�*z,�? %`t���_-� 1���E0�b8eO?a?�4gnpURGE_E�NB3��v�u�WFF�0DO�v��vWi���4�q*�WRUP_�DELAY ��CΡ5R_HOT �%�f�q:�.O�5R_NORMALH�
�OrOAGSEMI�QOwO�OlqQSKI%P-3���>3x$�O  _1_C_]&ot_b_ �_�_�_�_�_�_�_o (o:o o^oLo�o�o�o lo�o�o�o $�o H6X~��h� ������D�2��h�z�����$RB�TIF�4G�RCV�TMOU\��]���DCR-3��I� �QE=�U4�1D͛�C��JA?͜6��ט]���q��6��1�B�AY�����_V�R_ ;��x5;��0;��i;�du;�?t�<!��h��R���̝����� &�8�J�\�n�����������RDIO_T?YPE  4=���¯EFPOS1 ;1�C�
 x/:� H2��b�M���/��E� οi�˿ϟ�(�ÿL� �pς��/�i��ϵ� �ω�߭�6���3�l� ߐ�+ߴ�O����߅� ����2��V���z�� ��9����o����� ��@�R�����9���������OS2 1��;+�u���-��Q<���3 1������G���gS4 1�~���Z�E~�S5 1� %7q��/�S6 1Ũ���/�/o/�/&/S7 1�=/O/a/�/??|=?�/S8 1��/��/�/0?�?�?�?P?SMASK 1�߯� )�OF�7XNO�ܯFUO_C�MO�TE���X4uA_CFG �|M�1\A��PL_RANG�xA���AOWER ����@�FSM�_DRYPRG �%�%y?!_�ET?ART ��N/ZUME_PRO�O�_�_X4_EXEC_ENB  ����GSPDdP�P�X����VTDB�_�ZR�M�_�XIA_OPOTIONφ�����pAINGVERS6.a�z_�)�I_AIRPURƿ@ @O�o�=MT�_�0T�@zO��O�BOT_ISOLEC=N�F�1�a�e/NAMERl�bo�:�OB_ORD_N_UM ?�H�a�H721 � V1wLqr��qrV0qr�sps�u\@��PC�_TIMĖ��xު�S232�B1�����aLTEA�CH PENDA1N΀�7\H��x?�c�Mainte�nance CoKnsV2�#�"��_�No Use ��N��r���������С�rNPO>P�r\A�<e�qCH_LfgP�|Nw�	<�~�!UD1:b�z	�R�0VAILRq�2e��upASR + �:a�B��R_INTVAL�1f��I�+n��V�_DATA_GR�P 2���qs0DҐP�?`��?��o� �������կï��� ��-�/�A�w�e��� �������ѿ��� =�+�a�Oυ�sϕϗ� ���������'��K� 9�[߁�oߥߓ��߷� ���������G�5�k� Y��}��������� ���1��U�C�e�g� y��������������	+Q?uDA�$�SAF_DO_PULS�pE@�C�N� CAN�r1f�v�pSC�@�'��'Ƙ�QWV0D�DP�qL�L�+AV2 y� '9K]o��������ڈJ��2($Md($�C!u�1#
) @��Co/�/�/�.W)k/ �M��$�_ @݃T:`�/??&?~39T D��3? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO�|O֏��i%��O�O�O܉�!L� �;W�o݄�p�M�
�t��Di�pp�L��J� � ��jL���j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:����/c�u��������� Ϗ��B�%�1�C� U�g�y���������Ƒ��0RMS�EW]� $�6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬϾ����� M���*�<�N�`�r� �ߖߨ��������� �&�8�J�\�ǟ���� ������������� �,�>�P�b�p����� ����������% 7I[m��� ����!3EWit�OB3t �����//// A/S/e/w/�/�/�/�/��/�*��/?6���\R?�M	�12345678�XRh!B!S̺���� �?�?�?�?�?�?�?O OA�>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_o]-O�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�oq_BH�o�o�o! 3EWi{���������v[;�j�A�S�e�w��� ������я�����`+�=�O�a�xYD�k� ������ɟ۟���� #�5�G�Y�k�}����� ��v_ׯ�����1� C�U�g�y��������� ӿ���	�ȯ-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�� �ߕߧ߹�������� �%�7�I�[�m����v6�����z��!�3�O:Cz�  A�z   ��@�2�v0�� @�
���  	�r��������,����ph�u�����K]o��� �����#5 GYk}��0� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-?G��������*@  <X4t��$�SCR_GRP �1�'� '�� t �t�� E5	 ��1� �2�2�4��W1G3�;97�7�?�?OC���|�BD�` D���3NGK)R�-2000iC/�165F 567�890��E���RC65 �@��
1234�E�6Dt�A�����C�1�F�1�3�1)�1A�:�1�I	��?_Q_c_�u_�_���H��0 T�7�2�_�?@�_�_o�6�t��_@Lo�_poB8boK�h�@��UO��  u�P�1BǙ�B��  B�33B� �`�e�b�c�1Ag��oG  @t��e�1@>@�	  ?�w�bH�`2�j�1F@ F�`\rd[o�s �������*� �9�a�a)rU�@�R�d�v�B����ʏ��� ُ����H�3�l�W� ��{���Ě2C�?���7���9�t�!q@"p>SԪD_�U��r�`y��`ȏ�@�G�L�3��ϯ�A>G��1��"oe��)�t� �<�N�\�*��q�}���^� P���(����ӿ�g1E�L_DEFAUL�T  �D���t���HO�TSTR� ��M�IPOWERFL�  K����?�W�FDO� S�R�VENT 1�����P0� L!�DUM_EIP�翬��j!AF�_INE��ϵ!'FT�������9!�_B� ��i��!RPC_MAINj�LغXߵ�|�'VIS��Kٻ���o!TP��PU����d��M�!
PM�ON_PROXYN��e<���g���f����!RDMO_SRV���g��1�!R�DM���h, �}�!
~�M����il���!RLScYN�@����8��>!ROS��<��4a!
CE>�MTCOMb���kP�!	vCO�NS���l��!}vWASRC ����m�E!vUSBF��n4�0� �����/�'/��K//o/�RVI�CE_KL ?%��� (%SVCPRG1v/�*�%2�/�/� 3�/�/� 4??� 56?;?� 6^?c?� 7�?�?� H\��?L19�?�;�$ H�O�!�/+O�!�/SO �! ?{O�!(?�O�!P? �O�!x?�O�!�?_�! �?C_�!�?k_�!O�_ �!AO�_�!iO�_�!�O o�!�O3o�!�O[o�! 	_�o�!1_�o�!Y_�o �!�_�o�!�_{/�"�  �/� F�E1��� �����
�C�U� @�y�d���������� Џ����?�*�c�N� ��r��������̟� �)��M�8�_���n� ����˯���گ�%� �I�4�m�X���|������ǿ�ֿρ*_D�EV ���oMC:�H'�?GRP 2ׇ�+p�� bx 	�/ 
 ,y�ϒ� +r~ϻϢ�������� ��9� �]�o�Vߓ�z� ���߰������#�z� G���k�}�d����� ����������U� <�y�`���������*� ��	��-QcJ �n����� �;"_FX� �������/� /I/0/m/T/�/�/�/ �/�/�/�/�/!??E? W?�{?2?�?�?�?�? �?�?O�?/OOSO:O LO�OpO�O�O�O�O�O _^?�O=_�Oa_H_�_ �_~_�_�_�_�_�_o �_9oKo2oooVo�ozo �o�o _�o�o�o#
 G.@}d��� �����1��U� <�y����o��f�ӏ� ̏	���-�?�&�c�J� ��n��������ȟ� ���;���0�q�(��� |���˯���֯�%� �I�0�m��f������ǿ������R�d ��	�4��X�C�|�gϠϯ�%�����R������������ ���+��O�=�s߁� �Ϧ���i��������� �	��Q��x��A� �����������Y� �P���)���q����� ������1�U���I ��Ym���	 �-�!E3U {i����� �//A///Q/w/� �/�g/�/�/�/�/? ?=?/d?v?-?O?)? �?�?�?�?�?OW?<O {?OoO]OO�O�O�O �O�O/O_SO�OG_5_ k_Y_{_}_�_�__�_ +_�_ooCo1ogoUo wo�_�_�oo�o�o�o 	?-c�o��o S�O����� ;�}b��+������� ��ɏ�ݏ�U�:�y� �m�[��������ş �-��Q�۟E�3�i� W���{����دꯡ� ï���A�/�e�S��� ˯���y��ѿ��� �=�+�aϣ���ǿQ� �ϩ����������9� {�`ߟ�)ߓ߁߷ߥ� ������A�g�8�w�� k�Y��}������ ��=���1���A�g�U� ��y����������	 ��-=cQ��� ���w���) 9_���O� ���/�%/gL/ ^//7///�/�/�/ �/�/?/$?c/�/W?E? g?i?{?�?�?�??�? ;?�?/OOSOAOcOeO wO�O�?�OO�O_�O +__O_=___�O�O�_ �O�_�_�_o�_'oo Ko�_ro�_;o�o7o�o �o�o�o�o#eoJ�o }k����� �="�a�U�C�y� g�������ӏ���9� Ï-��Q�?�u�c��� ۏ��ҟ�������)� �M�;�q�����ןa� ˯��ۯݯ�%��I� ��p���9�����ǿ�� ׿ٿ�!�c�Hχ�� {�iϟύ��ϱ���)� O� �_���S�A�w�e� �߉߿����%߯�� ��)�O�=�s�a���� ���߇�������%� K�9�o������_��� ��������!G�� n��7����� �O4F�� g�����'/ K�?/-/O/Q/c/�/ �/�/��/#/�/?? ;?)?K?M?_?�?�/�? �/�?�?�?OO7O%O GO�?�?�O�?mO�O�O �O�O_�O3_uOZ_�O #_�__�_�_�_�_�_ oM_2oq_�_eoSo�o wo�o�o�o�o%o
Io �o=+aO�s� ��o�!���9� '�]�K��������q� ��m�ۏ���5�#�Y� ������I�����ßş ן���1�s�X���!� ��y���������ӯ	� K�0�o���c�Q���u� �������7��G�� ;�)�_�Mσ�qϧ�� ��ϗ�ߓ��7�%� [�I���Ϧ���o��� �������3�!�W�� ~��G��������� ��	�/�q�V������ w�����������7� .����O�s� ���3�' 79K�o��� ���#//3/5/ G/}/��/�m/�/�/ �/�/??/?�/�/|? �/U?�?�?�?�?�?�? O]?BO�?OuOO�O �O�O�O�O�O5O_YO �OM_;_q___�_�_�_ �__�_1_�_%ooIo 7omo[o}o�o�_�o	o �o�o�o!E3i �o��Y{U�� ���A��h��1� �������������� [�@��	�s�a����� �������3��W�� K�9�o�]��������� ��/�ɯ#��G�5� k�Y���ѯ������ {�����C�1�gϩ� ��ͿW��ϯ������� �	�?߁�fߥ�/ߙ� �߽߫��������Y� >�}��q�_���� ������������� 7�m�[���������� �����!3i W������}�� �/e�� �U����/� /m�d/�=/�/�/ �/�/�/�/?E/*?i/ �/]?�/m?�?�?�?�? �??OA?�?5O#OYO GOiO�O}O�O�?�OO �O_�O1__U_C_e_ �_�O�_�O{_�_�_	o �_-ooQo�_xo�oAo co=o�o�o�o�o) koP�o�q�� ����C(�g� [�I��m�������ُ � �?�ɏ3�!�W�E� {�i�����؟��� ���/��S�A�w��� ��ݟg�ѯc����� +��O���v���?��� ��Ϳ��ݿ��'�i� Nύ�ρ�oϥϓ��� ������A�&�e���Y� G�}�kߡߏ������ �ߵ��߱��U�C�y��g���������$�SERV_MAI�L  ���~��OUTPUT����RV 2�؍�  � (����_���SAVE����TOP10 �2�9� d  	��������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/�}/�/�/�/���YP�|���FZN_CF�G ڍ����j��!GRP� 2��'&� ,�B   A=0��D�;� B>0� � B4��RB{21l�HELL�"C܍�$�L�M�7|�?�;%RSR�? �?�?O�?%OOIO4O mOXOjO�O�O�O�O�O��O_!_3^�  �R3_a_s_AR_� ��{_�R�P)�xWIR2��d�\�]|�Rh6HK 1�v; �_o"ooFo oojo|o�o�o�o�o�o �o�oGBTf~b<OMM �v?��g2FTOV_E�NB��A�$��ROW_REG_UI����IMIOFWD�L�pߥ~@5�WAIT�r�Y�8��r�v@�0�TIM�u7��j�VA��A�>�_UNIT�s��v$�LC�pTRY�w�$���MON_�ALIAS ?e�yH�he��%�7� I�[�i�������� m����
��.�ٟR� d�v�����E���Я� �����*�<�N�`�� q�������̿w��� �&�8��\�nπϒ� ��O���������߻� 4�F�X�j�ߎߠ߲� ���߁�����0�B� ��f�x����Y��� ��������>�P�b� t�������������� (:L��p� ���c��  �6HZl~)� �����/ /2/ D/V//z/�/�/�/[/ �/�/�/
??�/@?R? d?v?�?3?�?�?�?�? �?�?O*O<ONO`OO �O�O�O�OeO�O�O_ _&_�OJ_\_n_�_�_ =_�_�_�_�_�_�_"o 4oFoXooio�o�o�o �ooo�o�o0�o Tfx��G�� ����,�>�P�b� ���������Ώy�����(�:���$S�MON_DEFP�RO ����c� �*SYSTEM�*M�RECALL� ?}c� ( ��}tpcon�n 0 >192�.168.56.�1:7188 8� .*=��11620 ԑ۟�����}7copy f�rs:order�fil.dat �virt:\tm?pback\Ü���Z�l�~��.#�mdb:*.*8���R�������2x#�:1\��-���8 ֯g�(y����3#�a+�=� ��W������1��� կf�xϊϝ�8���S� ����������Q�b� t߆ߙ���<�Ͽ�������
xyzra?te 11 ���ߠ��c�u���0��:�pickup.tp��emp�ϼ�U������
��/��lace��J���e�w����#�61?�U�B� T�����	������ cu�����>P� �*��_q ���:L��/ &��[/m//� �6/H/�/�/�/�/"/ �/�/�/i?{?�?�/2?�D?V?�?�?O�?��360�?�?cOuO�O��tpdisc 0-O0 ?OQO�O�O _Ƣ��O�O�Oi_{_ �_��1�1MT_�_�_	o �.��_R_couo�o� ,ϵ�Hi�o�o�o�Ϥ� �o7G�ocu�߭� ?�;CV����߯ �>@�h�z����o�o :U���
���A ӏd�v����,�@�� �����+���O�`� r���?)A-�?�Q������O+N3700 ��ӯd�v����_�_ >�<�T����	�o.o�� ӿd�vψϛ��� 6�I��������$����ʸ��d�v߈ߚ��$�SNPX_ASG 2������� >P��%�����  ?����PARAM ����� ��	��P�������*����OFT�_KB_CFG � �ô՞�OPI�N_SIM  
��%��������RVQSTP_DSBk�%�����SR �� �� &��ONRO�D��0���TOP�_ON_ERR � /�W�L�PTN� ����AH�RING_�PRMV� ��V�CNT_GP 2q��'��x 	�������� ��$��V}D��RP 1���(���_q� ������ %7I[m��� �����/!/3/ Z/W/i/{/�/�/�/�/ �/�/�/ ??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_r_o_�_�_ �_�_�_�_�_�_o8o 5oGoYoko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c� ����������Ϗ�� ��)�P�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ܯٯ����!�3��=PRG_COUNTL���[�_�'ENB��Z�M��N����_UPD 1�>�T  
H��� ۿ���(�#�5�G�p� k�}Ϗϸϳ����� � ����H�C�U�gߐ� �ߝ߯��������� � �-�?�h�c�u��� �����������@� ;�M�_����������� ������%7` [m����� ��83EW� {������/ ////X/S/e/w/�/ �/�/�/�/�/�/?0?�+?=?O?x?s?�?Q�_INFO 1�ɹ�� �F��?�?�?�O�9�]MEA??�>>�O�7���PA6��SB��u��P�YSDEBUG�i�ʰ�0d��z@S�P_PASSi��B?�KLOG ��ɵ���0�>H�?  ����1?UD1:\�D�>�B_MPC�Mɵ:_$L_ɱ�Aj_ ɱV?SAV ��MA��A�B�5 XSV�nKTEM_TIM�E 1��G��S 0���4�lXl_��0��T1SVGU�NSİj�'����`ASK_OPT�IONi�ɵ�����?a_DI�@��[eB�C2_GRP 2��ɹ�U�o�0@� � C��cP��`CF�G �k�\ �V�f`
EOB -Rxc���� �����>�)�b� M���q���������ˏ ��(��L�7�p��� �Vn���n�ϟ�\��� ��;�&�_�q^�Qd T�������ѯ����� ��)�+�=�s�a��� ������߿Ϳ��� 9�'�]�Kρ�oϑϓ� �����Ȭ�����1� C���g�U�wߝߋ��� ���߳�	���-��Q� ?�a�c�u������ ������'�M�;�q� _��������������� 7��Oa� �!�����! 3EiW�{� ����/�/// S/A/w/e/�/�/�/�/ �/�/�/??)?+?=? s?a?�?M�?�?�?�? O�?'OO7O]OKO�O �O�OsO�O�O�O�O_ �O!_#_5_k_Y_�_}_ �_�_�_�_�_o�_1o oUoCoyogo�o�o�o �o�o�o�?!?Q c�o�u���� ���)��M�;�q� _�������ˏ���ݏ ��7�%�G�m�[��� �����ٟǟ���� 3�!�W�o������� ïA��կ����A� S�e�3���w�����ѿ ������+��O�=� s�aϗυϧ��ϻ��� ����9�'�I�K�]� �߁߷�m�������� #��G�5�W�}�k�� ������������1� �A�C�U���y����� ��������-Q ?uc����� ����/A_q ������/�� �$TBCS�G_GRP 2���� � �  
 ?�  J/\/F/�/ j/�/�/�/�/�/�/;�#"*#�1,d0�?1?!	 H�D 6s33�[2�\5O1B�x!x?�9D)�6�L�ͣ1>����g6�0CF�?�?�8fff�1�>��!OI/Cj��6�1H4?B�C{OO�)H��0|A�]0@HD�O_O)H�1�8CFr�O�M@ �. XU&_ �O_Q_n_9_K_�_�_��[?��0�Sp �	V3.00�R�	rc65�S	*`�T"o�V|A��0 8 `�Y �G`mHo  � ��%@�_�o�c#!J2�*#�1-�o�hCFoG ��;!,C!�j�B"]b�l|�BPz� Pva����� ����<�'�`�K� ��o�������ޏɏ� �&��J�5�n�Y�k� ����ȟ������\ 	��-�ן`�K�p��� ������ޯɯ��&� 8��\�G���k����� !/ۿ�����5� #�Y�G�}�kϡϏϱ� ����������C�1� S�U�gߝߋ��߯��� ��	����?�-�c�Q� ���Y����m���� ��)��M�;�q�_��� ��������������% I[m9�� �����!E 3iW�{��� ��/�///?/A/ S/�/w/�/�/�/�/�/ �/?+?��C?U?g?? �?�?�?�?�?�?�?O O9OKO]OoO-O�O�O �O�O�O�O�O_�O!_ G_5_k_Y_�_}_�_�_ �_�_�_o�_1ooUo Coyogo�o�o�o�o�o �o�o	+-?u c����y?�� ��;�)�_�M���q� ������ݏ����� 7�%�[�I�������� o�ٟǟ����3�!� W�E�{�i��������� ï�����A�/�e� S�u����������ѿ �����+�a��y� �ϝ�G��ϻ������ '��K�9�o߁ߓߥ� c��߷�������#�5� G���}�k����� ����������C�1� g�U���y��������� ��	��-Q?a �u����� ��/���q_� ������/%/ 7/�/m/[/�//�/ �/�/�/�/?�/?!? 3?i?W?�?{?�?�?�? �?�?O�?/OOSOAO wOeO�O�O�O�O�O�O �O__=_+_M_s_a_ �_C�_�_}_�_�_ o9o'o]oKo�ooo�o �o�o�o�o�o�o #Yk}�I�� �������U� C�y�g���������я ����	�?�-�c�Q� s�u��������ϟ� �)�;��_S�e�w�!� ����˯��ۯݯ�%� �I�[�m��=�����pǿ���վ  ��� �)����$TBJOP_G�RP 2�ݵ��  ?���	A�H��O���� ���pXd�� ���� �� �,� �@�`�	 �D� ��CaD����`���ff=f��>��H�ϻ��L��	�<!a����>���=�B�  Bp��8�C��D)�U�CQp߃D�S�Ι�q�y���v� ?�������\<����U����%�CV�+��/���S�D5�mi�{Բ��ع�<����z�>�\>�33C� � CA��`�K�j���u�bߐ���z�;�9bB�E��>�׵ҳ� C�V���s����&���ǌ��;��6���%�]�D&� C��������
Ѷ�� ?s33����<wZ;u���ff���K������U�) C-_i�u�� ����*I@cM������������	V3.�00f�rc65e�* e��/ '� F�  F��� F� F��  G� G�X G'� G�;� GR� G�j` G�� G��| G� G��� G�8 G��� G�< H�� H� H���2 Ez  E��@ E�� E�B F� FR FZ F��� F� F��P<"G � G�pL#?h GV�� GnH G��� G�� G��( =u=�+�(�$`Q��?2�3?��  ��M?[:A���*SYSTEM�
!V8.3021�8 �38/1/2�017 A y�  p7M�TP�_THR_TAB�LE   $ �$�1ENB���$DI_NO���$DO�4  ���1CFG_T � 0�0MAX_IO_SCAN�2wMIN�2_TI�2DME\��0@�0�  � $�COMMENT �$CVAL�	CT�0PT_ID�X��EBL�0NUMQBENDIJfAZI�TID]B $DUMMY13���$PS_OVE�RFLOW�$��F�0FLA�0Y�PE�2�BNC$GLB_TM�7�EF@��1�0ORQCTR�L�1�$DE7BUG�CRP�@2@�  $SBR�_PAM21_V�P T$SV_ERR_MODU�4SCL�@RACT�IO�2�0GL_V�IEW�0 4w $PA$YtR�ZtRWSPtR�A�$CA@A�1�u_SUeU �0�N�P3@$GIF63@}$eQ lP_S��PiQ LpP�VI�<P�PF�RE�VNE�ARPLAN�A�$F	iDISTA�NCb��JOG�_RADiQ@$JOINTSPy��TMSETiQ�  �WE�UAC�ONS2@B�RON�FiQ	� $�MOU1A`�$LOCK_FOL�A��2BGLV@CGL��hTEST_XM�@@raEMPE`,Rx�b�B`�$US;A�fPH`2P�S�aN�bMP_�`�aQ�CENEdRr $�KARE�@M�3T�PDRAhP;t2aV�ECLE�32dIU��aqHE�`TOcOLH`�0qsVI{s{RESpIS32�y;64�3ACHX`�`�~qONLE�D29��B�pI�1  �@$RAIL_B�OXEHaPRO�BO�d?�QHOWWAR�0�r�@�qOROLM�B�A�C� �SK�r�@�0O_F9�!��S�qiQ�
>o �RVpOC:iQ_�SLOGaK�Y.a`ROUZbR��eAELECT�E<P`�$PIP�fNODE�r�r�q�IN�q2^��pCO�RDED�`�`}�S�0P9P@  wD �@OBAU`TA�a����C�@��p�P�q0��ADRAܥ0F@TCHup 7 ,�0EN�2�1A�a_�Tl�Z@�B�ObVWVA!A� � ApeR�5P�REV_RT�1�$EDIT��VS�HWR9�S@	UАI�S`yQ$IND�0@1QB蓗q$HEAD�5@ ��p5@溒KEyQ�@CPS�PD�JMP�L��5�0RACE�4U�a�It0S�?CHANNEzp��	WTICK{s�1M�`A�0@�HN�A�D0^�]D�`CG�P8���v�0STYf��q�LO�A�3B���jP� t 
��Gr�%�$���T=PS�!$UNIGa5A�E��0�FPORT��SCQU5ptR���B��TERCJ@*b�T=SG� �PPL6�$�DE��$`Thqb�0OK@>CV�IZ�D4�Q�E�APR�A�Ͳ�1��PU}aݵ_�DObk�XSV`KN�6AXI��7�qgUR_s�E$T�p���*��0FREQ_,hp<�ET=�P�b�OPARA`@.P
@�:[���ATHr�3@a�D�s�s�0 �2�SR_Q�0l8}��@�1TRQIc���$`�@��BRup��VyE@@��NOLD��AAp7a��x@�A��AV_MG����¨/���/�D)�D;�D�M�J_ACC.�C��<�CM��0CYC0M@3@��M@_E������٘@NbSSC��@  hPD1S���1�@SP�0*�AT:����@��i��B�ADDRES{sB���SHIF}b�a_W2CH�@&�I�@�|��TV�bI�2�]��h>��C�
�j
⎂V����0 \��������웱�@��CnӞ�aºꯆ:R����TXSCREE���0�TIN!AWS�P;��T��>�>�jP TQ�7P�B �6QP��
��
�>��RROR_"a�@����E�UEG�# ���U��@SXQ��RSM�� �UNEaXg��6��0S_�S���	0��>�Cx�b��o� 26�UE���2GRU�ͰGMTN_FL�Q�#POHgBB�L_�pWg@�0 �����O�Q�L1En���pTO`C��RIGH�BRD<ITd�CKGRg@��TEX,���WIDTH�sݐB�A�AZ{q��I_/@H���  8 $�LT_ �|�Y0@R�yP�b�s�w�B��GO�u��0D0TW� U�� �R�b�LUM8�!�^�ERV��]P�FP`>��1'@^r�GEUR�cF\���Q)��LP�Z�Ed��)'�$(�$(T�p#)5!+6!+7!+8"b�>CȰ`��Fj�q�aS�@E�USReT  <ġ�/@U�R��RFO�Chq�PPRIz�mx�@?A� TRIP�q�m�UN�0�4!�P ��0�5�7��b;�5� "T� ̱G �T7���}�&O2OSNAd6RA���;3wq�1#n_�S�^�2H���P�bU!"A$�?�?+"��;3OFFT�` P%O��3O@� 1#PD,D$NPGUN#K`S�B_SUBBPk 'SRT�0��&��"a�vp��OR�p�ERA�U���DT�Ib��VsCC��H�' ��C36MFB1���PPG?�( �(b`�STE�Q0ʀ9PWTѠPE����GXd) ����JM�OVE��{Q6RAN�4`?[�3DV�S6RLIM_X�3qV�3qV\X vQk\:V1�IP�2VF��C砽@��2G�*��IB�P
,�S� _�`�p�b��^�@ (0GB��� "P�@��pr+Gx �r �,�t�Rn@��s C@TeD#RI�PSfQV!�wd�Ԑ��D�$MY_UBY�$\d�;QA�S����h�q�bP_Sh�ף�bL�BMkQ�$j�DEYg�E�X� ���BUM_M�U6�X�D<q US��?��;VGo�PACI�TP�<Uyr�3`yrkSyr:;qREn�r�1l�8dyr�@,^�BTARGPP��q8eR{0�@- d���;cB	:r��RF�DSWqp�Sn�:s˰O�!d�Av�3���EE��U�p0m��v+HK�.��K�AQ0��0���?SEA�����WOR�@3��uMR�CVr/ ��O*��M�@C�	ÂC�sÂREF��̆ ��gRj�
�� Ȋ�ي���=�̆r�_RC ��s�����@����bp���:bo0 �Т��;��� �e�OAU���r��\c(`+�u���2��<���̰� �-=���f�K�SU�L3a.�C7Po/+p�NT�a��]���ag��g��!g�&�L��c���c������!R�@T��s�1���>o@AP_HUR�ۥ�SA>SCMP��FP�����_&�R�TP������X.��Q�GFS�E2d ��M� � Y0UF�_�����J��RO`� ����W,rUR�#GR�mq�I���D_V_h[D�@zY��3�WIN.rH���X-�V
A�RqR�P�W Ew�w�q|c6v,q��RvLOiPtc�PMc���3t +=�PA�' =�CACH 6����ŵ�,p����K�jۓC�QIo�FR"�qT� $֭�$HO�@�R��`�rc��[�`֘p��ڔ�VP�r<����_SZ3p���6����12� ��]pآ؆P��WA3�MP\��aIMGx����AD�qIMRE�ٔ6�_SIZ�P���!po�6vASYN�BUF6vVRTD�h�t�F�OLE_C2D�T��t��0C0a�Us��QP�X�EC;CU�xVEM�p��<��#�VIRC��VTP�����G�p���t��LA�s�!���QMco4��;�C/KLASQC	��ђ�@5  �A�� �@&B�T$��$`��6� |F@o���Xñ�T@�o�?a��"�uI��جr/��`BG� VEJ�`PK|p1���֖��0��HO+��R7 � }F���E�SLOW}w]RO>SACCE*@-�=�xVR:��11�yrcAD�/0rPA�ԩ&�D�1�M_qBa�81��JMP����A8y�b�$SS�C6u��M��C��@9$2��S8��N/�PwLEX��: T��C�Q��6�FLD6?1DEZ�FIQ r�O�qty��BVP2>��;� ϱP�V多�MV_PI Z��G�BP��`а�FIQ�PZ�$��������GA�%p�LOO0Tp�JCBT*����� ��ړPLAN�R&�L��F���cDV�'M �p���U�$�S�P.q �%�!�%#�㱶C4rG����RKE�1�VANC]G�A.0p <�@�?�?R_A�a = �?q??T0�9� Q3�@G> hܰ�	��K9��fA2b<X@̠OU�e�ݒA��
O���SuK(�M�VIE�p2= S0:�|R�? <{@XMԊ`U�MMY����Reڟ�D����1CU��`b�U�@@ $��@TIT 1$�PR8�UOPT?�VSHIFʀ�A`�a���T�0l����$�_R$�UړQ.qZ�U�s�o�t�Qav�Q5fST�G@cVSCO��vQCNT���3� }w�RlW �RzV�R�W�R�XLo^oTpjjA2��51D>a��0� �pSMEO��B%X�J�@�1u���_���@C4%�Gi�LI� ��^'��XVR�DDY��@T�� ZABC�P�E�r�bM��
.�1ZIP�EF%��KLV��L����b�MPCF�eGy��$p?�rDMY_LN$@Ar8��d�H ���g��>�M�CMİC��CAR�T_Xq�P�1 O$JvsptD��|r�r�w���u���U�XW�puUXEUL�x�q�u�t�u�q��q�y�q�v��Z�e�I Hk�d���Y��`D�� J 8xo�	V�EIGH�ƭH?("��f��9
�ĔK �= �C,���`$B&�K���1�_�B��LgRV� F8^���COVC؀qr@fq9��@}�e�
��4��7�D�TRȰ?�9V�1�SPH� Ǒ�L !�S�i�{� ����ST�S  �������0�`�0u�<�ѐNa1 ��w�� ����������������������"��	���a������*���������1N��RDI������@ğ֟����t�O|����������ίஔ�Sz��� >�����ſ׿ �����1�C�U�g� yϋϝϯ��������� �v�}���8�!�3�E� W���'�9�K�]���l� ����U�5` �0�0����0��@A�v�^`BF_TT��ի����I�V>0�2J�_��I�R 1&� C8����%к� ��C�  ��������� ���"�4�F�X�j�|� ������������1 gBTjx�����р���8�0B QI�Z lJ������� ��/"/4/F/X/F� ��t/�/b*���/�/��ԋbv�@`�v�MI__CHANU� `� #3�dV�`�u�&0�ET>�AD ?*��y0�m��/�/��?�?�d0RLPs��!&�!�4�?�<SNMASKn8��1_255.4E0�3�3OEOWO�OOLO�FS^Q �`�$X9O�RQCTRL �&�V�m��O��T �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo(l�OKo:ooo��;PE�pTAIL8�J�PGL_CONF�IG 	����/cell/�$CID$/grp1so�o�o1�#��?\n��� �E����"�4� �X�j�|�������A� S������0�B�я f�x���������O�� ����,�>�͟ߟt�@��������ίB�}c� ��(�:�L�^���`o��e��b���Ϳ߿� ��\�9�K�]�oρ� ��"Ϸ���������� #߲�G�Y�k�}ߏߡ� 0������������ C�U�g�y����>� ������	��-���Q� c�u�������:����� ��);��_q ����H�� %7�[m����]`�U�ser View� �i}}1234?567890�
/ /./@/R/Z$� �cz/���2�W�/�/��/�/??u/�/�3 �/d?v?�?�?�?�??�?�.4S?O*O<ONO `OrO�?�O�.5O�O �O�O__&_�OG_�.6�O�_�_�_�_�_�_9_�_�.7o_4oFoXo@jo|o�o�_�o�.8#o �o�o0B�oc�ir lCamera��o�@�����NE� ,�>�P��j�|�������ď�I  �v�)� �&�8�J�\�n���� �����ڟ����"�4�[��vR9˟���� ����ȯگ�����"� m�F�X�j�|�����G� Y�I7�����"�4� F��j�|ώ�ٿ���� ������߳�Y����� Z�l�~ߐߢߴ�[��� ����G� �2�D�V�h� z�!߃unY������� ������B�T�f��� ��������������Y� "i{�0BTfx� 1����� ,>P��Y��i�� ������/,/ >/�b/t/�/�/�/�/cu9H/�/?!?3? E?W?�h?�?�?F/�?��?�?�?OO/O�j	�u0�?jO|O�O�O�O �Ok?�O�O_�?0_B_ T_f_x_�_1OCO�p�{ ._�_�_oo+o=o�O aoso�o�_�o�o�o�o �o�_�u���oOa s���Po��� <�'�9�K�]�o� PEc����͏ߏ�� ��9�K�]������� ����ɟ۟����ϻr� '�9�K�]�o���(��� ��ɯ�����#�5� G��;�ޯ������ ɿۿ���#�5π� Y�k�}Ϗϡϳ�Z��� ��J����#�5�G�Y�  �}ߏߡ����������������   ��N�`�r��������������   $�,�J�\�n����� ������������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/�t/�/�  
��(�  �B�( 	 �/�/�/�/�/? ?8?&?H?J?\?�?�?ж?�?�?�*4� �n�O1OCO��gOyO �O�O�O�O��O�O�O _VO3_E_W_i_{_�_ �O�_�_�__�_oo /oAoSo�_wo�o�o�_ �o�o�o�o`oro Oas�o���� ��8�'�9��]� o����������ۏ� ��F�#�5�G�Y�k�}� ď֏��şן���� �1�C�U���y����� ���ӯ���	��b� ?�Q�c����������� Ͽ�(�:��)�;ς� _�qσϕϧϹ� ��� ���H�%�7�I�[�m� ��ϣߵ�������� �!�3�E�ߞ�{�� �������������� d�A�S�e�������� ������*�+r� Oas������0@ �������� ��)fr�h:\tpgl\�robots\r�2000ic6_�165f.xml �`r�����0��/����/3/ E/W/i/{/�/�/�/�/ �/�/�//
?/?A?S? e?w?�?�?�?�?�?�? �??O+O=OOOaOsO �O�O�O�O�O�O�OO _'_9_K_]_o_�_�_ �_�_�_�_�__�_#o 5oGoYoko}o�o�o�o �o�o�o o�o1C Ugy����� ��o��-�?�Q�c� u���������Ϗ��:K � 88�?�� 2��.�P�R�d����� �����П���(� R�<�^���r�����ܫ��$TPGL_O�UTPUT |���� ����%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ�Пϱ�����ˠ23�45678901 ��������0�8��� ��_�q߃ߕߧ߹�Q߀������%�7���} A�i�{����I�[� ������/�A���O� w���������W����� +=����s� ����e� '9K�Y��� ��as�/#/5/ G/Y/�g/�/�/�/�/ �/o/�/??1?C?U? �/�/�?�?�?�?�?�? }?�?O-O?OQOcO�? qO�O�O�O�O�OyO֡}�_)_;_M___q_]@��_�_� ( 	 ���_�_ o�_5o#oYoGoioko }o�o�o�o�o�o�o /UCyg�� ������	�?��Ƭ�-�G�u���c� ������ߏ���`�� ,�ΏP�b�@������ ��Οp�ޟ����:� L���p���$������� ܯ�X���$�Ư�Z� l�J������ƿؿz� ����2�DϮ�0�z� ��.ϰ��Ϡ�����b� �.���R�d�B�tߚ� �����߄����� <�N��r��&��� ������Z�l�&�8��� \�n�L���������� |����� FX�� |�0����� d0� fxV �����// �>/P/�</�/�/:/��/�/�/�/?
2�$�TPOFF_LI�M [��@W����A2N_SV�#0  �T5:P_MON S�S74�@�@2�U�1STRTCHK' S�56_=2�VTCOMPAT�J8�196VWVAR� j=�8N4 K�? O�@}2�1_DEFPR�OG %�:%?CONROD&O�?�_DISPLAY�*0�>?BINST_�MSK  �L �{JINUSER��?�DLCK�L�KQUICKMEN�OށDSCREP�S��2tpsc@�D�A1P6Y52GP_KY�ST�:59RACE?_CFG �Fr1��4.0	D
?���XHNL 2"�93��Q�; $B�_ �_o o2oDoVohozj��UITEM 2��[ �%$12�34567890<�o�e  =<�o�o<�os  !{!@�oZC�o{�o ���9K�o /��?�e����� �#���G���+��� O���ŏ׏Q�����͟ ߟC��g�y����]� �����������-��� Q��u�5�G���]�ϯ !����ſ)�տ��� q�ϕ�����3�ݿ�� ����%���I�[�m��� 	ߣ�c�u��ρ���� ��3���W��)��?� ���ߌ��ߧ����� c�S�e�w������ k��������+�=�O� ��s�EW��c�� ����9�o ��n���� �#�G�"/}=/ �M/s/�/��/// 1/�/U/?'?9?�/]? �/�/�/i?�??�?�? Q?�?u?�?PO�?kO�? �O�OO�O)O;O_�T�S�R�_UJ� 3 �bUJ �Q`_UI
 m_�_z_�_~8ZUD1:\�\���QR_GRP� 1�k� 	 @`@o!ko@Ao/oeoSo�own��` �o�j�a�_�o�o�e?�  '9{#Y G}k����� ����C�1�g�U�w���	�E��ÏS�SCB 2%[ �!�3�E�W��i�{�����\V_C�ONFIG �%]�Q]_�_���OUTPUT %Y�����S�e� w���������ѯ��� ��+�_A@�S�e�w� ��������ѿ���� �+�<�O�a�sυϗ� �ϻ���������'� 8�K�]�o߁ߓߥ߷� ���������#�5�F� Y�k�}�������� ������1�B�U�g� y��������������� 	->�Qcu� ������ );L_q��� ����//%/7/ H[/m//�/�/�/�/ �/�/�/?!?3?D/W? i?{?�?�?�?�?�?�? �?OO/OAOݟ�>� O�O�O�O�O�O�O�O _!_3_E_W_J?{_�_ �_�_�_�_�_�_oo /oAoSod_wo�o�o�o �o�o�o�o+= Oaro����� ����'�9�K�]� n��������ɏۏ� ���#�5�G�Y�j�}� ������şן���� �1�C�U�g�x����� ����ӯ���	��-� ?�Q�c�t��������� Ͽ����)�;�M� _�p��ϕϧϹ����� ����%�7�I�[�m� ~ϑߣߵ��������߀�!�3�E�W�i�LH�������s� ��hO������1�C� U�g�y���������t� ����	-?Qc u�������� );M_q� ������// %/7/I/[/m//�/�/ �/�/��/�/?!?3? E?W?i?{?�?�?�?�? �?�/�?OO/OAOSO eOwO�O�O�O�O�O�? �O__+_=_O_a_s_ �_�_�_�_�_�O�_o o'o9oKo]ooo�o�o �o�o�o�o�_�o# 5GYk}��� ���o���1�C� U�g�y���������ӏ����$TX_SCREEN 1������}��&�8�J�\�n���������ҟ��� ������P�b�t��� ����!�ίE���� (�:�L�ïp�篔��� ��ʿܿ�e�w�$�6� H�Z�l�~�������� ������� ߗ�D߻� h�zߌߞ߰���9�K� ��
��.�@�R���v� �ߚ���������k����$UALRM_MSG ?��� ��zJ�\� �������������������/"SFw+�S�EV  �E���)�ECFG ���  ��u@�  A� �  B��t
  x�s�0BT fx�������GRP 2�; 0�v	 �/�+�I_BBL_N�OTE �
T��l�r���q� +"DEF�PRO5�%9� (%k�/�p�/�/�/ �/�/?�/%??6?[?�F??j?�?!,INU?SER  o-/��?I_MENHI�ST 18��  �(�  ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1�?`OrO�O�O��9 (O:M936MO�O �O__�B/_A_S_e_ w_�_�_*_�_�_�_�_ oo�_=oOoaoso�o �o&o�o�o�o�o '�oK]o��� 4�����#��< V""A�_�q������� ���ݏ���%�7� Ə[�m��������D� V�����!�3�E�ԟ i�{�������ïR�� ����/�A�Я�w� ��������ѿ`���� �+�=�O�:�L��ϗ� �ϻ��������'� 9�K�]��ρߓߥ߷� ������|��#�5�G� Y�k��ߏ������� ��x���1�C�U�g� y�������������� ��-?Qcu`� rϫ���� );M_q�� ����//�7/ I/[/m//�/ /�/�/ �/�/�/?�/3?E?W? i?{?�?�?.?�?�?�? �?OO�?AOSOeOwO �O�O���O�O�O_ _+_.OO_a_s_�_�_ �_8_J_�_�_oo'o 9o�_]ooo�o�o�o�o Fo�o�o�o#5�o �ok}����T ����1�C��g��y����������O���$UI_PANE�DATA 1������?  	�}ӏ�`,�>�P�b�t� )v� ��V��şן���� ���C�*�g�y�`��� ���������ޯ���?�Q�8�u�R�� �A������Ŀֿ� ���_�0ϣ�B�f�x� �ϜϮ���'������ ���>�%�b�I߆ߘ� ߼ߣ�������7���T�Y�k�}�� ������J����� 1�C�U���y���r��� ��������	��- QcJ�n��0� B��);M� q������� /h%//I/0/m// f/�/�/�/�/�/�/�/ !?3??W?���?�? �?�?�?�?:?OO� AOSOeOwO�O�OO�O �O�O�O�O_ _=_O_ 6_s_Z_�_�_�_�_�_ �_d?v?4O9oKo]ooo �o�o�_�o*O�o�o�o #5�oYkR� v������� 1�C�*�g�N�����o "oӏ���	��-��� Q��ou���������ϟ �H���)��M�_� F���j�������ݯį ����7�����m�� ������ǿ����p� !�3�E�W�i�{�⿟� �����ϼ������/� �S�:�w߉�p߭ߔ���D�V�}����-�?�Q�c�u�)	��� ����������� ��� D�+�h�O�a������� ��������@R�9v	�`�Z��$U�I_POSTYP�E  `�?� 	 ����QUICKME/N  ����� RESTORE� 1 `�?  �i�!S`N�m~� �����/%/7/ I/[/�/�/�/�/�/ r�/�/�/j/3?E?W? i?{??�?�?�?�?�? �?�?O/OAOSOeO? rO�O�OO�O�O�O_ _�O=_O_a_s_�_(_ �_�_�_�_�_�O�_o "o�_Fooo�o�o�o�o Zo�o�o�o#�oG Yk}�:o��� 2���1�C��g� y���������d�����	��-��SCRE�� ?�uw1scHu2h�U3h�4h�5h�6h��7h�8h��USE�RJ�O�a�TI�j�k�sr�є4є5є6�є7є8ё� ND�O_CFG !����Ѩ PDAT�E ���?None _� ���_INFO 1"2`�]�0%3�x� 	�f�����˯ݯ��� ���7��[�m�P���ࣿ��ǿ�J�OFF�SET %� ԿσA֏�*�<�N� {�rτϱϨϺ�Ͼ� ���A�8�J�w�n� �ߒ�����
�����UFRAME � ʄ�G�RTOL_ABRT&��>�ENBG�8�G�RP 1&<?Cz  A���� ��������������:�� Ug��V�MSK  j�]�X�%N#���]�%�߫���VCCM�'����RG��*�	���ʄƉD � �BH)�p<2C�2)��PN?�` ��MR��20��p����"�р	 ���~?XC56 *�������N�5р��A@<C� ���ʈ)@;h�c���Rр|�Ђ B����6� t/T1/ /U/@/y/ d/�/�/�/�/*/�/	?��/???�c?u?��TCC��1��f�9��рр��GFSv�22w Й��2345678901�?�2ʈ"�6��?�!Oс>,12�QO_GB�@R 8N:�o=L����� ������OOA�O�O @O_dOvO�O�O�O�_ �O�O�___�_<_N_ `_r_Soeo�_Ro�o�_��_oo&o8o��4S�ELECF�j��$�VIRTSYNC� ��6�Bq�SIONTMOU4-tр��cu���3U��U��(�� FR:�\es\+�A\�o �� MC�v�LOG�   7UD1�vEX�с�' B@ ���qDES�KTOP-8U37T7F�6��q:�^��σ �  =�	 1- n?6  -��ʆ��xf,p�#�0=�̩ʹ���r�xTRAIN��2�1.���
. d��sq4w (,1��0�� )�;�M�_�q������� ��˟ݟ���I���crSTAT 5���@�o����E:$���ۯ�_GE��6nw�`. �
���. 2�HOMIN���7U��UC� �r�a�a�aCG��um�JMPER�R 28w
  ʯE:��suTs���� �߿���'�9�OϠ]ώρϓ�_v_�pR�E��9t���LEXr��:wA1-e��VMPHASE � RuCCb��OcFFLpc�<vP2�t�;4�04��8����b@�� �bb>?Gs33��Á�1�рL��ҕԈ�|��t�>x��Â�xf�o.���8/?P�X� $�2� x����0� ��� 6�+���l��\�j�|� ��������� �D� V���ZTf���� ������. �, BPb����� ��//(/:/� y/�b/��/�/L/ ? ??<?n/c?�/�/ �?�?�/�?6?�?�?�? OX?j?\O�?�OJO�? fO�O�O�O�O0O%_TO _xOm_�O�O�O�_�_ �_�__o>_P_EoWo �_xo�_�o�o�o�o���TD_FILTE:t�?�� ��Wp��]o$6HZl ~������ ��)�;�M�_�q�������SHIFTM�ENU 1@x�<��%����я�� 0���f�=�O���s� ����䟻�͟����P�'�	LIVE�/SNAPD�v�sfliv�b��{�ION G�yU���menu�����:�����±���A���	����b�K�S�5M����m`@�е���A�pB8��B����Ӝѝ�������m`� ;ӥ�/�M�E��uY��M�ֱ�MO��B���z���WAITDINEND�3���sOKN�.�OUT#�r�Sa�4�TIM�����GϮ�@π��`ϱ�ϱʞ�2�R?ELEASE���f�TM�����_ACTx��Ȫ�2��_DATA C��ի�%i��ߪ���R�DIS�b��$�XVR2�D��$�ZABC_GRPW 1E8�n`,@h�2��ǽZIP1�F�D� cCo������x�M�PCF_G 1G�8�n`0<o ���=�Hx8����t� 	�>w�  8R���0��e�����?�k�� ����5��
\�>�  �a � ����7������I��z��YLINuD�aJ�� �f ,(  *s��K�p���� �//+.mN/� r/Y/k/�/��/�/�/ 3/?�/�/J?1?n?U?`�/�?�?v�C�2K8��� ��O`o��7O~[Ol�?�Og���AA�ASPHE_RE 2LS�? �OX?�O__>_�?�O t_�_?�_I_/_�_�_ o�_]_:oLo�_�_�o �_�o�o�o�o#o l$7�ZZ� �k�