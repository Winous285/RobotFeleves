��   u��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����UI_CONF�IG_T  �� A$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]2�ODE�
3CWFOCA �4C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"��%�!BA�!j ?Ɵ"BG�%�!jIN=SR$IO}7�PM�X_PKT��"IHELP� M{ER�BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� GTB9I�:J�; &�USTOM0 �t $} RT_OSPID�,DC4Dn*PAG� ?^�DEVICEPIS�CREuEF���IGN�@$FLA�G�@C�1  �h 	$PWD_ACCES� E ��8��C�!�%)�$LABE� $Tz j�@�3�B��	CUSRVI| 1  < `��B*�B��APRIƍm� t1RPTR�IP�"m�$$C�LA�@ ��)�sQ��R��RhP\ �SI�qW�  �
�QIR�Ts1q_�P'2 L3�hL3!p�R	 �,��?�����Q�P�R�T�Q��R���P� � �T/o��
 ��zQQocouo�o�o�o�o Mo�o�o* <�o`r���� I����&�8�J� �n���������ȏW� ����"�4�F�Տj� |�������ğ֟e��� ��0�B�T��x��� ������үa������,�>�P�b��P/TPTX��򨅿ܗ��P sm����$/softpa�rt/genli�nk?help=�/md/tpmenu.dgd���� "�4��X�j�|ώϠ� ��A���������0� ��A�f�xߊߜ߮��� O�������,�>����zQ'`V�	bbS� ($�ߕ������������zQ�Q�c������*k
$m�d���
e�� c ��P����@�"*dn���	b�#`  �V������S�B 1�XR �\ }%`�REG VED��� whol�emod.htm�4	singlE�doub\t�riptbrows�@�!�� ��/AS|��/Adev.EsJl�o�1�	t���w�G/ Y/k/5/�/�/�/�/�/ ?� �P?*?<? N?`?r?�?�?�?�?�6 �@?�?�?�? O2ODO E	�/�/wO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_� �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-??z� ������
�� O@�R�!�3�����QO cOI�ݏ��*�%� 7�I�r�m�������� ǟٟ�����_/�)� W�i�{�������ïկ �����/�A�S�e� w�����iֿ���� �0�B�T�f�x�s��� ��}Ϗ����ϭ����� >�9�K�]߆߁ߓߥ� ����������#�5� ^�Y�k�9������� ��������1�C�U� g�y������������� ��ſ2DVhz� �������
� �@R	���� �����/*/%/ 7/I/r/m//�/�/�/ �/���/�/?!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSO! �O�O�O�O�O�O�O_ _0_+T_f_5_G_�_��_�Z�$UI_T�OPMENU 1��P�QR� 
d�QfA)�*defaul�tqOZM*le�vel0 *\K	G o� So�_�Qocbtpio[2�3]�(tpst[1�heo�ouo3oEo��-
h58E01�.gif�(	m�enu5&ypHq1!3&zGr%zEt4M{4�a������� ��eB�C�U�g�y������,�prim�=Hqpage,1422,1��ݏ� ��%�0�I�[�m��葟��2���class,5�����h�)�4���130�@f�x�������5���53ʏ���� �2�
5���8ٯm���� ����4�ٿ����!�3�^I�P�Q�_k�m�]��a[ϕ�o�ftyx�m�o�amf[0�o���	��c[164�g.�59�h�a���&tC8$|Gr2uK} ��azmWw%{�ߩsK� ]�6�H�Z�l�~�ɿ���������𢡊��80$�?�Q�c�u�����̐2����������	 ��ʟ?Qcu� (T�������Ѥ1.�N`r�������ainedic����//���config=single&��wintpĀ /`/ r/�/�/]J�QV¤/�/ e�/�o�o??1?D? U?g?y?�?�/�?�?�? �?�?	OO-O?O�aO �O�O�O�O�O�O��_ _*_<_N_`_�O�_�_ �_�_�_�_m_�_o&o 8oJo\ono�_�o�o�o �o�o�o{o"4F Xj�o|���� ����0�B�T�f� x��������ҏ���MNS�,�wω¯����w���s��<�����¡�u�͔�V�|�F7 ��7����԰�Οp�����6��u7��� �����/�A��227쯃�������˿Z� l�����,�>�P�/!$13�ϛϭϿ� �ϐ�����+�=�O� ��s߅ߗߩ߻����� "���'�9�K�]�����6d��������,$۬74r��/�A��S�e��,����%	TPTX[209�����24����������18�������
����0P2���1_��E�tv����\�Q�u10�1=��ïqC:4$treeOviewA#�3�&dual=oU81,26,4� ���n����	/ /-/�Q/c/u/�/�/$�/ֺ;@b�3`r �?)?;?F/_?q?�?@�?�?�?�/�/\2�/t2��O1OCO�?��1�/E���O�O�O�y6XO��edit� zO�O_._@_׹?�� �OCL_�_�_�_~��_ �_G�o}o�CoUo goyo�o�o�o�o/o�o �o	-?Qdu ӥ������� I?2�D�V�h�z���� ��ԏ���
���� @�R�d�v�����)��� П�������<�N� `�r�����%���̯ޯ ���&���J�\�n� ������3�ȿڿ��� �"��_�_X�o|��o ��ϱ���������� ߋ�)�S�e�x߉ߛ� �߿��ߓ��,�>� P�b�t￿������ ������(�:�L�^� p��������������  ��$6HZl~ �������  2DVhz� �����
/�./ @/R/d/v/�/7�IϾ/ m��/I���??)?;? M?`?q?�?�/�?�?�? �?�?OO%O7O��nO �O�O�O�O�O�O%/�O _"_4_F_X_�O|_�_ �_�_�_�_e_�_oo 0oBoTofo�_�o�o�o �o�o�oso,> Pb�o����� ����(�:�L�^� p��������ʏ܏� �/�/$��/H��?MOk� }�������ş؟�W� ���1�C�U�h�y��� ��_Oԯ���
��.� y�@�d�v��������� M������*�<�˿ `�rτϖϨϺ�I��� ����&�8�J���n� �ߒߤ߶���W����� �"�4�F���X�|�� �������e������0�B�T���*d?efaulta�2��*level8����������{� �tpst[1]���ytpi�o[23��u�������	menu7.gif�M
�13�	�5�
h��
�4�u6�
 ʯ?Qcu���� ����//�;/�M/_/q/�/�/�/6"�prim=�page,74,1�/@�/�/??+?6"�&�class,13 0?f?x?�?�?�?=?O25�?�?�?O O2O5#D<�?lO~O�O�O�O�/�"18�/�O__'_9_DON26@_u_�_�_�_�_��$UI�_USERVIE�W 1���R 
�A��_>��_
o�m(o Qocouo�o�o<o�o�o �o�o�o);M_ qo~���� ��%��I�[�m�� ����F�Ǐُ���� ��.�@���{����� ��ßf������/� ҟS�e�w�����F�P� ��̯>���+�=�O� a����������Ϳp� ���'�9��F�X� j�ܿ�Ϸ������ϐ� �#�5�G�Y�k�ߏ� �߳����߂������ z�C�U�g�y��.�� ����������-�?� Q�c���������� ����)��M_ q��8���� �� 2�m ���X���/ !/3/�W/i/{/�/�/ J�/�/�/B/??/? A?S?�/w?�?�?�?�? b?�?�?OO+O�/�? JO\O�?�O�O�O�O�O �O�O_'_9_K_]_ _ �_�_�_�_�_lX