��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�   � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d PPINFwOEQ/ ��L A �!�%/� H� �&�)EQUIP 2� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CES0s!_81F3K2> ��! � $�SOFT�T_I�Dk2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5Xk2S�CREEN_(4n_2SIGE0_?|q;�0PK_FI� �	$THKY�GPANE�4 ~� DUMMY1d�DDd!OE4LA!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTc@�D5�F6�F7�F8�F9�G0�G�GJA �E�GbA�E�G1�G ��F�G1�G2�B!S�BN_CF>"
 }8F CNV_J� �; �"�!_CMNT��$FLAGS<]�CHEC�8 �� ELLSETU�P � $H�O30IO�0� %��SMACRO�RR'EPR�X� D+�0��R{�T UTO�BACKU��0 �)DEV�IC�CTI*0��� �0�#�`B�S$�INTERVAL�O#ISP_UNI�O`_DO>f7ui�FR_F�0AIN��1���1c�C_�WAkda�jOFFu_O0N�DEL�h�L� ?aA�a1b?19a�`C?��P�1bE��#sATB�d���MO� �cE D [M�c���^qREV�BIL�rw!XI� QrR o � OD�P~�q$NO^PAM�Wp�t�r/"��w� �u�q�r�0D~`S p E �RD_E�pCq$�FSSBn&$CH�KBD_SE^eA�G G�"$SL�OT_��2=�� V��d�%��3RO��a_EDIm  � � �"���PS�`(4%$EP<�1�1$OP�0�2��a�p_OK�UST1P_C� ��dx��U �PLACI4!��Q�4�( raCOsMM� ,0$D冀���0�`��EOWB BIGALLOW�G (K�"(2�0VARa��@�2aI��L�0OUy� ,�Kvay��PS�`�0M�_O]����C�F�t X� GR�P0��M=qNFL�I�ܓ�0UIRE��$g"� SWIT{CHړAX_N�P]Ss"CF_�G�� �� WARN�M�`#!�!�qPLI��I�NST� CO�R-0bFLTR^C�TRAT�PTE�>� $ACC1a��N ��r$ORIأo"��RT�P_S�Fg CHG�0I���rTא�1�I���T�I1��� x i#�Q��HDRBJ; C,�U2'�3'�4'�5'�U6'�7'�8'�9s!:ҢO`T <F П�����#92��LLE�Cy�"MULTI�b�"N��1�!���0�T_}R  4F STY�"�R`�=l�)2`�����`T |� �&$c�Z`d�pb��P�MO�0��TTOӰ�Ew�EXT����ÁB���"�2� ��[0]�}R���b�}� D"}����Q����Q�kcG�� �^ȇ1��ÂM���P��� ŋ� L�  ���P��`=A��$JOBn�/��i�G�TRIG�  d�p�߻���³��7�����!CO_�M�b! t�pF̝ CNG AiBA � ����M���!���p � �q��0��P[`��,i�*�"6���0t�B񉠎"J��_Rz�gC�J��$�?�Jk�D�%C_�;������0ФR�t#�C ������G����0NHANC̳$LGa��B^a��� �D��A�`��gzRɡ�!��p�3DB�RA�sAZ�0KELT��\���PFCT&��1F�0�P��SM��cI��1�% ��% ��@R��a���� S��&���M 00{o Ve#HK~�A^S��h�����I_T$�"�6SW�CSXC�)�?!%��p)3��T�$@��PANN�&�AIMG_HE�IGHCr�WIDLI AVT�0��H F_ASPװ��`�EXP�1���CWUST�U��&��
|E\�%�C1NV q_�`�a��' \%1y�`OR�c,"�0gsdk��PO��LBSYI�G��aR%�`좔Psp�m��0G3DBPXW�ORK��(��$SKP_�`}��!<q�TRp ) ����P���� �0�DJ!d/�_CN��R�#� �'PL�S�Q�d�"s�DKA7WAw'����^A�@NFZpfBDBdU��*�"!PRS��7�
ЖQ����+ �[pr�$1�$-ZϢ�Li9,v?�3�ʠ��-�?�4C��.��?�4ENEy��� c/�?�3J0RE`���20H��CuR7+$L,C,$i3
��? =KINE@�K!_D�I�RO�`��祀��ȳqvC��h �FPiAÃ3uR�PRN�B��MR��U!�u�C�R[@EWM �SIGN��A� .q��E�Q-$P��g.$Pp 2�/ PB7�PT2�PDu`�L���VDBAR@�GO_AW���Jp �� �DCS�pZ�C�Y_ 1���@1�<�Q?fIG2�Z2>fN>�����
�qS&c~}P2 P $��SRB?�e�P=hPwgF�QBYl�`gT+1^�THNDG�23���KS�SE|�Q��SB!L㸣cc�TG1sQ=L�4 HpZ <���VTOFB�l�FEfA�ǿb�TqSW�5�bDOC���MCS�f�`Z$r�b �H� W0��T#�eS�LAV�16�rINP��f��LyqQP�_7� $,�S����=��v��uFI��r줭sc�!���!W1ԭrNTV�'��rV	��uSKIvTE�@W���:�&J_� _�00��SAFE�A�_S}V��EXCLU��*B �PDJ L1�k��Y�d�ƻrI_V<� !PPLY 0b�旁DE~w��_ML�2�B $VRFYi_�#��Mk�IOU@��憻 0���:�O�PƜ�LS�@jb;�35H72��Sr�� Px%�X�{P�hs� �� 8 @� TA� qঠ� �c_SGN��96����@�A� ����iPt!��s"��~UN�0jdՔ�U���B �@� ��� ����G1l�OGI.�2: @�`Fؒ���OT�@@�:41(��774C2�M`NIB�2;�R������A�qDAY1#LOA�D�T/4~�;30� �[EF�XI�b< @�%1O㠈3� _�RTRQ��= D��`@��Q@  B�EjP"�㥎�<��B�� 	�@��AMP��]>�a�����a�8Sq�DU�@q��.�"CAB��?A��0�NSs���IDI�W�RK�^�� V�WV�_]���> �D�I��q�@� /^.�L_SE2�T� ��/�Z`��0��#�CE_��u�v�j��SWJ�j� 𲰂�	�2��=c�OH�z�3PPJ�v�IR!��B� ��w�d��B"����BASh��� X ���V����?C��Q���RQDW��MS����AX}�8�u�LIFE� �7�A1CҁNJ���S��H���Chs�>��C`QaN"�U��OV� �_�HE����SUP$�hbC�� _�Ԥ�B��_����[Q��Z��W���ו�Tb��cXZ$ `1��Y2F�ECM@T��t@�N�p��G1��9A `��P.�HE��SI�Zy֥�u��BN�pU7FFI���p� ��Q/40�<26C3��M�SW9B 8�K�EYIMAG�CTM@A��A�Jr|#>��OCVIET���'C C�V L�t���s?� 	G1� :�D�"pST�!x�0�� 0��Ѡ��|0���EMAIL���@�� �ba_FA�UL��EH�CC�OU�p}$T@��F�< $���eS�]���ITvBUF@��q���T  ���	BdC�t����#��SAVb$)�e� �A� }���Pi�e@U�b`_ H���	#OT{BH�lcPր(0�
{��AX1#��� @��_GJ�f1YSN_�� Gj�D�UT/0e��M����T8�F��ِ�A!H�(@u���C_r@�@K�D�����=pR���uD�SP �uPC�I�Mb��J���U`��ЁEƀ��IP�sdu��D� �TH0ȸc��TuA�HS{DI�ABSC�ts��0Vzp*} �$,�#��NVW�G�#�$H0� FJ�/d�j�ASC��U��MER��uFBC3MP��tETH�!AmI��FU��DU 0�a�@;⠂CD�O �� ���R_NOA�UTg` J�`�Pp2��n4ĥPSm5�CF }5CI�.� �`k3� =KH *}1Lp��Q� �&�I���4#Q�6s���6ѡ�60��6���67
�98�99�:J��8�:U1J1J1J1+JU18J1EJ1RJ1_J�2mJ2�;J2J2�J2+J28J2EJ2�RJ2_J3mJ3�:3�KJ3J/�G8J3*EJ3RJ3_J4mB2q�EXT�>aLC` ��F�fF�5Q9g�5���FDR�MT��VC��C�wa}".C�REM,�FAj�OVM��eA�iT7ROV�iDTm �jMX�lIN�i���jN�IND�`!�
x<p /$DG�Ð�`opS�9�D��`R�IV)0Qbj�GEA-R�IO0�K�bu�Nj�x�.؎��p�q>j�Z_MCM>�C��d`��UR)2N ,<{1��? ��
 s?�pI�?�q�E���q0�T0lbO�����P� �RI�T5��UP2_ gP Ѡ#TD= @��C����qP�J�,�wBAC;Q T��h$9 O�)��OG���%E��3e&0IFI���e0�0����PT��6�FMR2ieRO vbY�vbLIq��{g���P�f��Ŗb_mAN~"F�_F�I4+�M;v`�r}DGCLF��D7GDY��LD�q>tA5[�5S�كk�S���M� T�FS� l�T P�)���|
�/$EX_)��@�)�1�� ��*�3�b�5b��G�!ieU� � p&2SWKO>��DEBUG�S���0�GRY�zU�#B�KU� O1�@ O�PO8��Π0l��ΠMS]�OO�V�SM]�Eq}��pQ`_E V �$�X����TER�M2�W;�6�ORI�Ā6�X;����SM�_��$7�Y;�XP�O�TAy�Z;�I�ON�UPB�[� -��QbV$|G���W$SEGź�אELTO��$wUSE0NFI�с��p���`���X$UFR����q0豘��D5h�OT1Ǵ TqA_ �C�NSTd��PATT!��Y�PTHJ!B0En�K0�ART� ���������REL��&S�HFTF"�_���_�SH��M�!B0x� ȃ�n���Z���OV9R
#&SHI�����U�2 �AYLO$ 5I1�_�d���d�ERV�0*�}  ��b?�d��Q�����A��RC
���AScYMh���WJ�apE�����f�2�U��d�5����D5��aP#Gи!	�ORd��M�h0GR!���\ ��΢�^�����Nk�] �E���TOC�졳q��OP��N z�3&1��e�aO�a> RE���R�#&O0��`�e��R]���������e$PWRSpIM���[�R_���VI1Sy�r���UD�t��� ^>�$H|����_ADDR9fH$�Ga�z�s�i1qR� =_ H8�S� ��S��C��C���CSE�abaHySO0��` $����_D`���P�R�aHT�T� UTH�a =({0OBJE1u𶎄$9fLEP�|-=b � *g.!AB_qT���Sk�#DBGLV�5#KRL"�HIT��BG0LO���TEM4$��b�������SS�p�4JQ�UERY_FLAD��f WYA���c��� PU�"B� 1��4G��H��H~B �IOLN~��d/0i�C��$�SL�� PUTM_�$���PwpܛrSLA�� e/2����ӡ����0IO F_AuS�f��$L�� U���#�04�#����,�HYOgN!'#؁� UOP�g `  l!9f�b>$�`E&�!��P����'�!E&�"��&�P_MEM�Bk0T h XF IPz�v��"_#0 v����0��Oc6�1�w�DSP�' $F�OCUSBGԃ�{UJhfi � 60�S��JOG�W2D[IS�J7��O�ү$J8�97��I�6!�2�77_LAB�Q����0�8�1APHMI�pQ�3�7D+��J7JRA4`P�_K�EYp �K^ILMON�j&`�$XR =0cWATCH_ �DӘ�&U1EL� �y`B&�k GpG�VP�-f�fBCTR��fB5� �LG|�l ���+h�"��LG_SIZ{Y��E
��F,
 �FFD�HI�H�H ��F�HM��F�@���C 5V
�5V
 5V�@5VM��5W�`S)@S���S��LNv1��mx �� ��R��4a�PÀU��Qk�L�S�RDAU�UEA I���R��PGH���� B�OO~�n� C-"2�ITGcd��)&�REC-jSCRN,)&DI(#S��RG����cl�!#��H�b�!Sa"Wkd�!�T!#JGM�gMgNCH"FN�2��fK�gPRG�iUqF�h	��hFWD�h�HL/ySTP�jV`�hĀ�h`�hRSgyH!�{&C�Es��!#���g�yUt�g �¬f|@6#�bG�i4�CPO�JzZeEsM�w�82�iEX'TUI�eIP�cw��c�� �c���`�a����s���Jg��KaNO{�ANqA"貇�VAI�0�zCL����DCS�_HI��������O�����SI)��S'��hIGN�@��C��aT����DEV��wLL��a_SBU𠔠oa@�mT��$�GEM'�9nD �EsAb�p�a@ЅC�!��O+S1��2��3��*83�����q �T0v�-�絡.e�IDX����-fL�b�STm R�PY0����� p$E��C ���  ����� ��r L*</��Q(06����6�EN 6��ՕKc_ s �Y��P$ dKaD� �{MC�Rt �T0�CLDPm ��TRQLI`��e0x�f��FL>1��_����DUA��LD������ORGe0�r���WX������Y���V�O�u � 	���uu���%Si�Tx��00�ް�S�[�RCLMC�i����{�m[�C0M9I��O�v d�Q6��RQ�00�DSTB��Y� ��{a���AX��@�� �EXWCES����M�
��wc �¹�������x(��_A@�ʊ l����V�K|��y \*�2��$M�BLIE��RE�QUIR����O���DEBU��L
�M{�zW�.!��B��i���N,03Ѩ�a{�R�RkHV�DCE�ƶTIN3 `!�TRSMw0p�S�N�����s�<�PST�  |nh�LOC9�RI� 9�EX��A��:���^��ODAQo%}��c$@�Q΂MF �A�_���p�C��P��SUP"� �F�X��IGG�"~ �0��MQ���v�5@� %����m ���m ����6#DATA����E� 1�NP" �N�� t�MD
IF)?�!��H���1!� �Q"ANSW�a!ܑS�
!D�)��H3Q�$�� ?�CU�@V0_ >0���LO�P$��=ұ���L2�p�����RR2I5��  ��QA�X� d$CALII��NUG�2g�RINp<$R�SW0��K�A�BC�D_J2SqE����_J3v
p1SP�@6 ��	Pp�3��\�����J���P�O村IM��[�CSKAP��$�P�$J�Q[�Q,6%%6%,'���_AZW��h!ELx�����OCMP�����1X0RT�Q�#�c1�c@�Y�1��(t�0�*Z�$SMG�p�����ERJ�N�IN� ACߒ��5�b��1
�_B�542d���414X҆>9DI~!�ãDH �30���c$Vo�Y�$�a$� ���Q�<�.A���ňH ��$BELy lH�A/CCEL?��8��>�0IRC_R��i���ATw�c�$P)S �k�Lm�yP D���0G�Q�FPACTH�9WG�3WG3&B��#�_�2�@�AV�r��C;@�0_MG|a�$DD�A@[b$FW(����3�E�3��2�HDE�KPPA�BN.GROTSPEE�B��_x�,!���DEFg��1m�$OUSE_��PzЉC ���YP�0V� �YN��A{`uV��8uQMOU�ANG��2�@OLGC�TINC~���B�D���W���ENCS���°A�2��@INk�I`&Be��Z�, VE�P<'b23_UI!<�^9cLOWL3��pc x��UYfD�p��Y�� ��Uy�C$0 fM3OS`���MO�����V�PERCH  vcOV�$ �g9��c ��\bYĄ��'�"_Ue@$0��A&BuLcT�����!ec�\jWvrfT3RK�%h�AY�s hчq&B�u�s���&l��Rx�MOM|���h� ﰞ ���C�sYC����0DU��BS_�BCKLSH_C &B��P�f�`}S�7���RB��Q.%CLAL���b?��pX�t�CH�Kx�H�S�PRTY�����e�����_�~��d_UMl�ĉC�у�ASCLބ PLMT�_L�#��H�E������E �H�-��Q#p_��hPC�a�hH��ЯE2ǅCw��XT�0�GCN_(N�þ���SF�1�iV_RG�e��!��&B���CATΎSH~�(�D�V᱀�f�'A�	� �@P�A΄�R_Pͅ�s_ y�뀎v�`x��s�����JG5�6Ф�G`OG|���rTORQUQP ��c�y�@�Ңb�q�@�_W�u�t�!�14�P�33��33�I;�II�I�3F�&������@VC�00���©��1��2�ÿ�¶�JR�K����綒 DBL�_SM�QO�Mm�_sDL�1O�GRV:�`3ĝ33ģ3�H_�8�Z@a�COSn˛ n�LN���˲��ĝ0 ��� ��e��ʽ̃��1Z���f�MY����z�TH��.�THE{T0beNK23�3�Xҗ3��CB]�CB�3C��AS���e�0�ѝ3��]�SB�3��Nh�GTS@! QC����'y��'����$DU��;w	��Q������qQ����$N	E$T�I�����)I7	${0L�AP�y��`�k�k�LPHn�W�1eW�S���������W���������{0V��V���0��V��V��V���V��V��V�V�H�����7������H��H��H��H��H�O��O��OTF	��O��O��O��UO��O��O�O�ƁFW�}��	�����S�PBALANCEl�{�LE��H_P�SP1��1��1��PFULC5\D�\��:1��!UT�O_��ĥT1T2��22N���2, �����q^<�-B#�qT�HpO~ �1$�INSsEG�2{aREV��{`aDIFquC91م('o21�dpOB!d�=��w2��7P��~�LCHWARR�2AB���u$MECH��ДQ�!��AX�qPB��&r�~2�� 
�"��1e7ROB�`CR r�%z��S0MSK_��4� P �_�OPR�1�2(47Qst1 �,`*R(0)cB�(0|!�IN!�MTC�OM_C���0� � �@0 �A$ONOREc�2�l �~2� 4�GR���%FLA!$?XYZ_DA��LP^;@DEBU�2 �0�lR�0� ($mQC;ODS� �2�r�� �p$BUFoINDX*PD�2�MOR3� H %0�p�0��:@�p�QB�"�1��NF�TA9Q0&@�r�G.B� � $SIMUL���0qxs�AsOBJE3>�FADJUS�H�@OAY_I��xD�G�OUTΠ�4�p�P_[FI�Q=8AT#� Y,`W�1P +�PQ�+ 9�uDjPFRI4 �PUT0�RO�
`�E+�Sp�OPWO���0�,@SY�SBUi� @$SO!P�QBy��ZU�[+ �PRUNn2�UPAB;0D�V�"�Q�`_�@F��PP!AB�!H��@/IMAGS�%0?��P!IMQAdIN�$��RcRGOVR!DEQ�R�@�QP�Pc�� L_��feÂ�ސRBߐ<pX�MOC_ED'@�  H��Ni M�bG��MYc19F�0EaSL3�0� x $OwVSL�SDIsPDEXǓ�f֓Hq�b	V+��eN�a
��Pp��cwx�bw��d_�SET�0� @0�Cr�%9�RI�A3�
Vv_��bw{qnq?q�-!�@� �4BT�� àATUS�$TRCA�@PB�s'BTM�w�qI�Q�d�4F��s�`0� DB%0E�P�b�rr�E1"�qQpd��qEXE��p���a�"��tKs��Rp&0�pUP�01�9$Q `XNN�w��x�d���y �PG|5�� $SU�B�q�%xq�q|sJM/PWAI$�Ps���LO ��1
 �E$�RCVFAIL_C@1�PÁR%P�0�#����Ȕ� �
�R_{PL|sDBTBá����PBWD��0UM��IG�Q `��,�TNL ��b�R eQ�2���qP��@�EǓ��֒��DEF�SP� � L�%0� ��_���CƓUCNI�S�wĐe�R)���+�_L
 P�q}0PH_PK�5���2RETRIE�|s�2�R���F�I�2� � $��@� 2��0D�BGLV�LOG�SIZ�C� ���Ud�"|�D?�g�_T:�ʥ!M�@C
 #EM⌭R��y0�8CHE�CKS�A��o01�B�0.�0R!�RNMGKET��@�3砹PV�1� h�`A�Rp� �1)P�2>�S��@OR|sFORM3AT�L�CO�`q�d���$Z��UX�P�!r?qPLIG�1��  ˣSWI�m �21AX,�G�AL_ � $�`@��B�a��CS2D��Q$E1��J�3DƸ� T�`P�DCK�`�!�RCO_J3����T1l׿� �˰C_Q��` � ��PcAY��S2u�_1|�2|�ȰJ3�Иˈ�x�Ɨ�tQTIA4��u5��6S2MOMK@@����������y0B׀�AD��������PU��NR��C���C����4�` I$PIN�u�41�ž� ��:q�R~ȇ��ٯ� �:�h��a�֬��ց��1�'1R\uSPEED G��0�؅�� 7浔؅�%P7�m�F�p�U��؅SAM �=G��7��؅MOV	B� e0�� ��c2 ��v��浐�� ���c2@nPsR����İ$QH���IN8�İ��?�[��6�؂A���X����G�AMM�q�4$GGET1R@�SDe�zmB
�LIBR[��y�I�7$HI�0_�5a@c2E`@#A@ 1LW^U�@	�1a¬&o�ʱC�=�n S`�p �I_��pPmDòv� ñ'����mD��	ȳ� �$�� �1��0IzpR� D`T#|"c���~ LE^1�41�qwa�?�|�M�SWFL�MȰSCRk�7�0��Ѻpv���Z 0�P�@�9@���2�cS_SAVE_Dkd%]�NOe�C�q^�f�  ��uϟ�}ɕQ��}��Ѐ}*m+��9��ժ(��D �@���������b3 1�RA�Qm�7
5�#���^��LVuԡ 7� �YL��
A
'�VAS	BtRna`7 GP�B
Bl3
A%`�$GSB1W? �2�2c�Ȭ3oBB1M&@�;CL �8���G�b�1v���9M!Lr� �N�X0�d$W @�ej@b �� @=�BD�BK�B �-�> �P����ycJİX �OL�ñZ�E����uԣ ��OM�R/d/v/�/��/��A�jM`��e�_��� |��H �� jV��yV��yP�ʗW�Vr��E��� IWJ������NTP=���PMpQU�� �� 8TpQCO�U,�QTHQ�H�OY2`HYSa�ES��aUE `"#�]O���   �P�0L�rUN�p�3��9O$�J0� P�p^e�������OGRA��qk22�O�d^eI�Tm�aB`INFOBI1���k�ak2���OI�b� (!SLEQ(��a��`�f�oaS� ��� 4�TpENABLBbpPTION|s����Yw\��1sGCF��O��$J�ñfb���R�x!�]ot�����_EDŀJ0� ��N��@K�᪃E�S NU�w�xAUT<,!�uCOPY����(�v�8 MN��^�PRUT�� ��N�pOU��$G�cbn���RGADJ�I1�2�X_B0ݒ�$ ����@��W��P������@㊀��EX��YCLB��NSr6u�N0�LGO��A�NYQ_FREQZ�W���+�p�\cLAm"����Ì�u�CRE  c� IFl�ѝcNA��%i��_GmSTATUxQPmMAIL��  1��yd����!���ELEM�� �|7 DxFEASIGq 2��v��q!�er$�  I�`�"��a�e�|I�ABUq�E�`D�V֑a�BAS��b� [�Ub�r % �$y���RMS_TRC�ñj���Cpa��ϑ�� ����C�YP	 � 2� g�DU�� ���Ԣ�0-�1��1����qDOU�ceNLrs��PR30;p�r�GRID�aUsBA�RS(�TYHs��O�TO�I1��P`_"��!ƀ��l�O�@7t�� � �`�@P�OR�cճ��ֲSReV��)���DI. T���!��+��+�U4)�5)�6)�7)�I8���F��:q�M`?$VALU|�%�� 0��7t�� !Cu'!�a���� (FgpAN#��R�p|0� 1TOTAL��,[��PW�It�&�REGEN$�9��S�X��sc0��Q���PT1R��Z�$�_S ��9дsV���t���rb�E��x�a�"^b�p��7V_H��DA�C�Ў��S_Y4!�B<�S��AR�@2� >f�IG_SEc��d�˕_b`��C_����w��?r��%�b�H�SLG#�I1��p@"=���4��S�2̔DE�U!Tf.p��TE�@����# !a����Jv�,"��IL_MK��z�н@TQ�P�a��T��2VF�CT�P���^�Mu�V1t�VU1��2��2��3��3��4��4����������1�"IN	VIB@N�; �!�B2>2J3>3
J4>4JI05����"���p�MC�_F`3 � LP!!�r�M= I���M� [PR��� KEEP_HNADD�!f�	C�A��!����"O�Q I����"���?�"REM9@!�ϲ^uzU���e!HPWD  �SBMSK"G�a	!B2B�
#?COLLAB�!@��2�����o��`�IT��A`��D�� ,pFLI@��O$SYN� ;,M�@�C>��%�UP_D�LYI1�MbDEL�Am ј�Y�PAD��A��QSKI�PE5� ��``O�n@NT�1� P_ ``�b�'�`�B]0�'�� �)3��)��)O��*\���*i��*v��*���*9��J2R‎���?sX��T%�|1��{2ܐ�|1�a���R�DC!F� ��pR"�sR�PM�'R^��:8b�2�RGE�p2��3d�FLG�Q�J�t��SPC�c�UM�_|0��2TH2N�P�F@o0 1�� �0EF�p11��� l[P�E-Ds#ATWo�[�w�B �`�d�A�p3�BfcA�HnP�B��_D2gB��mOO�O�O�O�O�G3gB��O�O_ _2_D_
�G4gB�g_y_�_�_(�_�_�G5gB��_�_�oo,o>o�G6gBŀaoso�o�o�o�o�G7gB��o�o&8
�G8gB�[m�H���ES����\@ǡ`CN�@�_@w-E��^� @o�L�m�IO�ፉI����^APOWE!� W�: �1���0�� �5%Ȃ$D�SB;���֒ �h C�L@��S232s�̓ ��0�u.��IgCEU{���PEV@>��PARIT�њ��OPB ��FLOW�TR2�҆]����CUN�M�UX�TA���INTEORFAC3�fU����CH�� �t� � ˠE�A$L����OM��A�0"נI���/�A�	TN���Tо ��ߓ��EFA� �"!�Ҏ��� u!��� �O�� &*�� ������  2� ��S�0�`�	�' �$3@}%:B��䎣�_���DSP���JOG��V�h�_P�!s�ONq0%�0����K��_MIR����w�MT7��A�P)�w�>@"���;AS�������;APG7�BRKH����G �µ!! ^���i���P���<����BSOC��w�N���16�SV�GDE_OP%�FSPD_OVR��u �DвӣOR$޷�pN��߶F_���6��OV��SF�<���
�F0����UF�RAF�TOd�LC1Hk"%�OVϴ ��W[ ���8�Ң��͠;�  @ BT�IN����$OFeS��CK��WD����������r���TRr��T�_FD�� �MB_C �B��B����(�.Ѻ�SVe��琄�}#��G)�<�AM��B_0��jթ�_M@�~�x�ቂ��T$CA�����De���HBKX�����IO�������PPA���������Տթ���DVC_DB��?����A���,�X� b��X�3�`���3�0����ϱU8󳠈�CAB�0��ˠ��c� �Ow�U�X��SUBCPU�ˠS�0�0�R�����!�A�R�ł�!$HW_Cg@A��!���F��!�p� � �$�U r�l�e�AT�TRI��y�ˠCY�C����CA���FLT ��������vALP׫CHK�o_SCT��F_e�cF_o����FS�J�j�CHA�1��98I�s�8RSD_!�0���恩�_Tg�7��� �i�EM,��0M"f�T&� @�&�#ޮDIAG��RAOILACN���M�0 �"��1���L���{�PRB�S   ��pC4�&�	��F�UNC�"��RI	N�0 "$�7h�� S_��(@��`�0p��`A��CBL� �u�A����D�Ap�a���LD@ܐð�����j���TI%��@�$CE_RIAAV��AF�P=�>#,��D%T2� C��a��;�OIp��DF_aLc�X��@�LML��FA��HRDYO,���RG�HZ 7�����%MULSE�� �����k$J�ۺJ����FAN?_ALMLV�1�WRN5HARD�r��Fk2$SHADOW|�A���O2 s�0N�r�J�_}����AU- R+�TO_SBR���3���:�e�6�?�3MPIN�F@{��4��3R3EG�N1DG�6C1V��s
�FLW��}m�DAL_NӀ:�����C	����a�vU�$�$Y_B�ґ u�_�z��7� �/�EGe����ð�AAR������2p�G�<�AXE��wROB��RED���WR��c�_�M��S�Y`��Ae�VSWWcRI���FE�STՀP����d��Eg�)�$�D-�{2��BUP��t\V��D��OTO�19)���ARY���R0���6�נFIE����$LINK�!GkTH�R�T_RS���E��QXYZt��Z5�VOFF��b�R�R�X�OB���,8d����9cF�I��Rg��􃻴,��_J$�F�貿S��q0kTu[6��1�w �ad�"�bCԀ+�DU�º�F7�TUR0X#�e�Q�2X$P�ЩgFL�Pd���@p�U�XZ8���� 1�J)�KʠM��F9�p��ӓORQ����fZW30�B�O Pd�,��t����A�t'OVE�q_BM���q ^C�udC�ujB�v�w0L�wg��tAN=�Q �qD!`A�q��=�}��q �u�q���dC��"���SERϡj	�E��HT�ńAs�@�Ue�X��W����AX ��F����N�R�� +��!+�� *�`*��`�*��`*�Rp*�xp*�1 �p*�� '�� 7�� G� � W�� g�� w�� ���� ��� ��đ��DEBU=�$8D3�h����RAB�����r�sV��<� 
�� i�`A��-񷧴���� ��a���a���a��Rq���xqJ$�`D"�R9cL�ABOb�u9�F�G�RO��b=<��B_���AT�I`�0`�����u���1��AND fp�ຄ���U���1ٷ ���0�Q�������PNT$0M�SE�RVE�y@� $�%`dAu�!9�PO��[0ЍP@�o@*��c�x@�  ]$]�TRQ�2
\�d�Bf��j�D"2�{��" � _ � l8"T�c6ERRub��I��VO`Z���TO	QY�V�L�@)�1R��J� G;�%�Q�2 [�T0e�� ,7�ř���]�RA#� 2'� d@����r�7 �Y@$�p��t ��OC�f���  ��COU�NTUQ�FZN_wCFGe�� 4B�F��Tf4;�~�\� ��
����uC� ���M: �"`A��U��q: �FA1 d�?&�X�@=����_B�A�<����AP��o@H�EL@���� 5�`B_BASN�3RSRF �C�Sg�!��1
ש�2���3��4��5��6���7��8
ל�ROaO�йP�PNLdA��cABH�� ��AC-K��INn�T��GB�$Uq0� +\�_P�U��@0��OUJ�P�HH���, u��T�PFWD_KAR���@��REGĨ P��P�]QUEJRAO�p�`2r>0o1I0������P����6�QSCEM��O��� A�7STYk�SO: �4DIw�E���r!�_TM7CMANR�Q��PEND�t�$KEYSWIT�CH���� HE��`BEATMW3PE�@LE��]|� �U��F>��S�D_O_HOMB O>�6_�EF��PR>a9B(�ABPx�CO�!��#�OV_M�b[0# �IOCM�d'eQ�ъ�HKxA� �D�QG��Ue2M������cFORC�CWAR�"�O}M�@ � @r�T:#�0UHSP�@1&U2&&3&&4�A�*s�O��L"�,�HOUNLO��c4j$�EDt1  �S�NPX_AS���� 0+@ @��W1$�SIZ�1$VA����MULTIP�L��#! A!� � $��� N$S`�BS�ӂAC���&OFRIF�n�S���)R� NF�ODBU$P���%B3=9GŸ�Ҫ�y@� x��S�I��TE3s�r�cSKGL�1T�R$p&���3a�P�0STMTd1q�3P�@5VBW�p��4SHOW�5���SV��_G��� Rp$PCi�oз��kFB�PHSP' 1Av�Eo@VD�0vC��� ���A00޴RB% ZG/ ZG9 �ZGC ZG5XI6XI7�XI8XI9XIAXIB�XI ZG3�[F8PZGFPXH��XdI1qI1~IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1 Y1Y1YU2WI2dI2qI2~I2�I2�I�`�X�IQpT�X�I2�I2�I2�I2 Y2Y2Y�p�h�dI3qI3~I3�I3��I3�I3�I3�I3��I3�I3�I3�I3� Y3Y3Y4WI4�dI4qI4~I4�I4��I4�I4�I4�I4��I4�I4�I4�I4� Y4Y4Y5�y5�dI5qI5~I5�I5��I5�I5�I5�I5��I5�I5�I5�I5� Y5Y5Y6�y6�dI6qI6~I6�I6��I6�I6�I6�I6��I6�I6�I6�I6� Y6Y6Y7�y7�dI7qI7~I7�I7��I7�I7�I7�I7��I7�I7�I7�I7� Y7Y7TF��0P� Uc�� l�נ��
>A820�����RCM2���MT�R��|���Q_��R-��ń�����[�YSL�1�� � �%^2��-4��'4��-Y�BVA�LU�Ձ���)���F�J�ID_L���H�I��I��LE_������$OE�S�Ab�� h �7�VE_BLCK�¡1'�D_CPU7ɩ 7ɝ ������E���R � � PW��>�E 6��LA�1Saѝ������RUN_FLG�Ŝ������ ����������H���Ч����TBC2��� � _ B��� b�r� W?�eTDC����X��3f�S�CTHe�����R>�~k�ESERVEX��e��3�2 �d���� �X -$��LENX��e����RA��3�LOWI_7�d�1��Ҵ2 �MO/�s%S80t�I���"�ޱH����]�DyEm�41LACE��2�CCr#"�_M�A� l��|��TCV����|�T�������0Bk�)A�|�)AJ$��%EM7���J��B@Rk�X�|���2p `�0:@q�j�x JK��VKX�����ы�J0����JJ��JJ��AAL���������4��5�Ӵ NA1�� ����LF�a_�1� ѡ �CF�"�� `�GROUP���1�AN6�C�#~\ REQUIR�Ҏ4EBU�#��8�$Tm�2���|�ё %�� \�A�PPR� CA�
�$OPEN�CLOS<�Sv��	k�
��&� �<�M�hЫ���v"/_MG�9CD@�C ���DBRKBNOL�DB�0RTMO_�7ӈr3J��P ��������������6��1�@ �	�$��� � ���'��-#PATH)'B!8#B!��>#� � �@�1S�CA���8INF��UCL�]1� C2@UM�(Y"��#�"������*���*��� PA�YLOA�J2L�ڠR_AN`�3L���9
1�)1CR_�F2LSHi2D4L�O4�!H7�#V7�#ACRL_�%�0�'��$��H���$H�C�2FLEX�:�J#�� P�4��F߭߿���0��� :����|�HG_D�����|���'�F1 _A�E�G6�H�Z�l�~����BE�������� ����*��X�T,�C� ���@�XK�]�o�^Av�	T&g�QX>�?��4T X���eoX�������� ����������	-	:�J@� �/�M0_q~�۠AT�F��6�ELHPѬs�Jڗ � JEoCTR�!�ATN���v|HAND_VB�q�1��$� $:`�F2Cx���SW�Ms��� $$M,00�_Y�n i��P\����A��� 3����<AM��_AmA|��NP�_UDmD|P\ G���E�STaM�nM�NDY��� C���� 0��>7_A>7Y1�'��d�@i`�P��������"Qs$�� O�4D'"��J����ASYMl%A��� l&��@�-Y1�/_ �}8� �$��� ��/�/�/�/3J	<�:p;�1�:9�D_VI��x���V_UN!I�ӝ��cF1J���� 䕶�Y<��p5Ǵ�y=�6��9��?�?>�wc|�4�3  �$� �ASS  ����s�=��|�h�V�ERSIONp����
��I�RTU<�qσ�AA�VM_WRK 2� �� �0  �5�z�������� �	8�)�L�=���!�:�w�^�|�(ܛ݀��7ѭ���������B�SPOS� 1���� < ��A�S�e�w���� ����������+�=� O�a�s����������� ����'9K] o������� �#5GYk} �������/�/1/C/U/ⰑAXgLMT��X#�%�7  dj$INs/�!�i$PRE_EXE��(� �&)0�q��������LARMRE?COV �ɥ"�
�LMDG �����[/LM_IF �ˆ!X/c? u?�?�?�:Q?�?�?�?< OM, 
0�8O��4�cOuO�O�O�NGTOL  ���A   �O�K��{PP)�O ; ?6_,_>_P_{� $BR_�_w�o_�_ �_�_�_�_o�_'oo7o]o�!��O�o�o�o �o�o�o�o+=�Oa�PPLIC�AT��?��� ��%@Han�dlingToo�l �u 
V8.30P/33�@�lt��
88�340�slu
�
F0�q�z=��
2026�tlu���_��7DC3�pJ  ޭsNonelx� �FRA�������B�TI�V�%�s�#��UT/OMOD� E�)�P_CHGAPO�N������ҀOUP�LED 1���� ��"�4�uz_�CUREQ 1���  � >�>��*ސ�4��!��x�=~� ��u���Hm����HTTHKY����w��� 7����%�C�I�[�m� �������ǯٯ3��� �!�?�E�W�i�{��� ����ÿտ/����� ;�A�S�e�wωϛϭ� ����+�����7�=� O�a�s߅ߗߩ߻��� '�����3�9�K�]� o�������#��� ���/�5�G�Y�k�}� ������������ +1CUgy�� ����	'- ?Qcu���� /��/#/)/;/M/ _/q/�/�/�/�/?�/ �/??%?7?I?[?m??��P�TO�@�����DO_CLEAN�܏��CNM  �K >�aOsO�O��O�OD�DSPDR3YRO̅HI��=M@NO_'_9_K_]_o_ �_�_�_�_�_�_�_J�MAX�p�4�1��뇂aX�4"��"���PLUGG���7���WPRC�@B;@?K_�_ebOjb�O��/SEGFӀK�o�g �a;OMO'9K]�o�aLAP�O~Ǔ �������/��A�S�e�w���΃TO�TAL-fVi΃USWENU�`�� ���䏺�P�RGDIS�PMMC�`{qCL�aa@@}r��O�@�f�e��_STR�ING 1	ˋ
_�MĀS���
`�_ITEM1j�  n������ ����Ο�����(� :�L�^�p����������ʯܯI/O �SIGNALd��Tryout �Modek�In�p�Simula�tedo�Out�.�OVERR~�@ = 100n��In cycl�"�o�Prog OAbor8�o���Statusm�	�Heartbea�ti�MH Fa�ul����Aler ���ݿ���%�7�pI�[�m�� �3 f��1x���������� �*�<�N�`�r߄ߖ� �ߺ����������WOR�`f�L���&� t����������� ��(�:�L�^�p���p��������POd� ����d���%7I [m����� ��!3EWi��DEV���� ����//'/9/ K/]/o/�/�/�/�/�/��/�/�/?PALT��81d�?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O&?GRI`f��AP? �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o@o$o6oHo�OR�� �a�OZo�o�o�o�o�o &8J\n��������noPREG<>%��o�L� ^�p���������ʏ܏ � ��$�6�H�Z�l��~�����$ARG�_L�D ?	����ӑ�  	$�W	[�]�����ƐSBN_CONFIG 
ӛ�&�%� �CII�_SAVE  ��E�<�ƐTCE�LLSETUP �Ӛ%  OM�E_IO��%MOV_H�������REP�l���UT_OBACKt�0�FRA:\�� ���_�'`r���=�� J� 	�������ͿĿֿ�6���� 	�1�C�U�g�yϋ�� Ϸ���������ߜ� 5�G�Y�k�}ߏߡ�,� �����������C�U�g�y����a��  )�_�_\A�TBCKCTL.�TMP DATE.D;<��	��-�?�.�INI;0p�8���MESSAG�T�^�_�ېi�ODE�_D��W�8�H���Ox����PAUS���!�ӛ ((O֒��
��*N <r`��������"����TSK  ��=�C�	��UPDT��\�d����XWZD_E�NB\�4��STAp[�ӑ�őXIS&�?UNT 2ӕ`�� � 	 ����0@��n��b{N�G�7���`�`9'$7�  /L/�^. "YK��ާď` �Ď}��=/�/pa/�/�/�MET�`2�P�/?�/<?��)SCRDCFG� 1C`��\�\�1?�?�?@�?�?�?�?6��QX� �??OQOcOuO�O�O O �O$O�O�O__)_;_0�O�O���GR��X��zS��NA��қs	�wV_EDZ��1e9� 
 ��%-��EDT-`h_ʪ�_o�`/A����-��_�	�������_�o  ���e2�oɫko�o�6k��o!hozo�o�c3 Y�o��o�n��4F�j�c4%��r� ��nN��� ����6��c5�a�>����n�@��̏ޏt���c6�� -�
�Q��n�Q�����@�Ο�c7����֯� �n���d�v�����ca8U��_����0
 }�~��0�B�ؿf��c9!ϑ�nϵ� }Jϵ�`��Ϥ�2φaCR�o į9�K����������n���zP�PNO_D�EL�_xRGE_U�NUSE�_vTIG�ALLOW 1��Y~�(*S�YSTEM* 3�	$SERV_G�R�R 69���REG�B�$d� <9�NU�Mg��z�PMU|�� 5LAY� � <PMPA�L[��CYC10�����������UL�SU��{�����D��L�N�BOXOR=Ik�CUR_;�z�PMCNV���;�10���T4�DLI�%9�[�� �ߨ��'9K�]oR�zPLAL_?OUT Dcc��QWD_ABOR���	��ITR_R�TN���Y� NO�NS8� �CE_RIA_I���<F_1���B =[_PA�RAMGP 1.�w`_�x���Cp  .U� � � � U� � � � U� � � � o�  D5`D$T3!g-�<$�H$�T$_� DX � eX "� B�D1� -9X @� 6?� <{HE��ONFIy����!G_P��1� �e�U??�0?B?T?f?x?�?�!KoPAUSX�1�UR ,Z��?�?�? �?�?OOOTO>OxO bO�O�O�O�O�O�O_�2O_ey�P�COLLECT_�_�Y5auGWEN���I�cR QNDE�OS�W���1234567890�W�S�u�_�VNy
 H�y)�_ #oS��_ohoT�AoSo �owo�o�o�o�o�o�o <+�Oas �������� \�'�9�K���o��VQ�2W[ � t�VIO �YcQy�H&�8�J�\��T-R�2؍(��1
��j��  �����%�_MOR҂!� + �'� 	 �5�#�Y�G�}�k�����Ӂ"��2? �!�!3 ҡ�Kڤ��$R_#*_	��>�C4  AS y�C  x�A3!z'  BC!�PB/!�P�C  @*��z��:d�
�UIPS$���T���FPROG % �*6߼�8��I�����&RҴKEY_TOBL  )VR�� �	
��� !"#$%&�'()*+,-.�/�W:;<=>?�@ABC��GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~��������������������������������������������������������������������������������͓���������������������������������耇�������������������s���1��LCKۼ83���STA�д�_AUT��O(��U�INDtTD�FQ�R_T1_�Q�T2`��7$����XC�� 2����P8
�SONY XC-�56�������@���u� ���А�HR5���cT0�B�7T�f�A�ffrꬿ����  �������5�G�"�k� }�X��������������ǼTRL��L�ETEG��T_�SCREEN ��*kcsc�:U$MMENU� 1&�)  <���y�� Ã�=&s J\������ �'/�/]/4/F/l/ �/|/�/�/�/�/?�/ �/ ?Y?0?B?�?f?x? �?�?�?�?O�?�?CO O,OyOPObO�O�O�O �O�O�O�O-___<_ u_L_^_�_�_�_�_�_ �_�_)o oo_o6oHo �olo~o�o�o�o�o �o�oI 2X�h�z���� _MANgUAL�ߕ�DB���L+�DBG_E7RRL��'��� �\�n���~�NUMLIMK��d �p�DBP�XWORK 1(�I�ޏ����&��ŽDBTB_@ �)��������qDB_AWAYz�_�GCP  ��=�װ�~�_AL��D�z��Y��M �� �_)� 1*����
͏�����6�@�_M{�IS�AЉ�@B�P�ONT�IMJ� ���p�ƙ
�ۓMOT�NEND߿ڔRECORD 10}�� �>�?�G�O����?���2�D�V� h���p������*�߿ �Ϛ���9Ϩ�]�̿ �ϓϥϷ�R���J��� n�#�5�G�Y���}��� �����������j�� ��C��g�y���� ��0���T�	��-�?� ��c���\�������� ��P�����;��_ q�����(�L %�4[� ����^t�l !/�E/W/i/{//�/ /�/2/�/�/??�/�z�TOLEREN�C��B�В��L����CSS_CNSTCY 116�'  ?Β�?�? �?�?�?�?�?OO&O 8OJO`OnO�O�O�O�O��O�Oc4DEVIC�E 126�  b�*_?_Q_c_u_�_�_��_�_�_�_?�d3HN�DGD 36��Cz�^LS 24]�__oqo�o�o�o�o�o�_e2PARAM 5�B��t�d�c4SLAVE �66�e_CFG� 7��gd�MC:\e0L%0?4d.CSV�o���c|�r�"A �sC	H�p&a&��n��
w��f�r���<�ÀJP�>��\�_CRC_OUT 8U����oEp?SGN 9U�Ƣ���\�16�-OCT-22 �14:21�p��02��4��9V? UBu1�݁��nހ��o��Im��P�uG���@uVERSION� ��V3�.5.11E�EF�LOGIC 1:^ݫ 	6���|�C���^�PROG_ENB����͢��ULS{� ��^�_ACCLIM|���Xs��WRSTJN[���ţ�^�MO��¡Zr,�INIT ;ݪ�s5� *�OPT�$p ?	i�B�
 	R575�cV��74��6��7��#50��R�Ƣ2��6���X�y�TO  Ѕ��?�Y�VP�DE�X�d���@W�P�ATH A��A�\E�����7;IA�G_GRP 2@��k,�"	 �E�  F?h Fx E?`�D��û��V1"�üb��T0K�9�Cf�p}y�pY�dC�pq�B�i�ù�mp4m5 �78901234�56��;���� � A�ffA��=qAةpх�A��HAĩp��������A���Mk���@��tpX�p��W0A�T0T0�pB4ü Qô����
���(�A�A�
=A�L����A��
A_�Q�A��������e�����e�� Pe�:��{A�Jd�����dѩp���_���A���������r߄ߖߨߺ߾@�EG�A@�p:��RA5d�/��)*��#P�d�l�������"�4�F�@�Pz��AJ��c�?��9�p�A3\)A,/��A&����0@��������@�cP�_]��AW�P�UJ��C��<d�4�-d�%G��(�:� L�^�@���$H Z��.|���� bt� 2Vh �xm�����[���s������=�
==��G��>�Ĝ���7���8�{�b�7�7�%��@ʏ\"&�pi�.%��@�Ah�p�9 A��<i���<xn;=R��=s��=x<��=�~Z�;���%<'�'�~ ��?+ƨC� � <(�U� �4"����&��!��%ùf��@?Œ ?�?@?R?g��$^? �?"?�?�?�?�?�?��?)7L?S�FNB$�/"Eͽ�>OG�ΐԬq���sD�L4�x�CA� �Gb�tφ���-_7_�C���_;�/_�NE�D  E�  EOh� D[PbRD_�¿�_�8�?��p(ج�Q��
'��Y�Q4����3�P������QħѪC=�/�D"	�q<�{_�_w_o�K:o@bù��Y7m�)6;��T*�/9B�Po�o
o�o�o�o��o�oĿDICT_�CONFIG ΂�Yt؃�eg��ԱSTB_F_TTS�
ę�Vs3���
�iv[�M�AU���Y�MSW�_CF*pB�  ��Q�OCVIEWf}pC�}���6� 
��.�@�R�d�w� ������ȏڏ�{�� "�4�F�X�j������� ��ğ֟������0� B�T�f�x�������� ү������,�>�P� b�t��������ο� �ϓ�(�:�L�^�p�,���|RC�sDJ�r!ϐκ��������7�&�[�otSBL_�FAULT E����xu�GPMSK�_w��pTDIAG� F.y�q�I�UD1: 67�89012345��;x�MP�o!�3�E� W�i�{��������������/�A��( W!�J�"
��v�TRECP����
 �����M�(: L^p����� �� $6]�o��l��UMP_OP�TION_p�ގT�R�r`s���PM�E^u�Y_TEM�P  È�33B�pp �A  ��UNI�pau!�vY�N_BRK G��y��EMGDI_�STA%�1!G%NmCS#1H�{ �K ��9�/_}dd�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO��O�O �O�O�I�!�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXo�JO�o�o�o�o �O�o�o+=O as������ ���'�9�K�]�wo ���������oۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�o�]������� ɏ�����	��-�?� Q�c�u���������Ͽ ����)�;�M�g� y��ϕϧ�]�ӯ���� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�_�q�{��� ������������/� A�S�e�w��������� ������+=O i�s������� �'9K]o �������� /#/5/G/ak/}/�/ �/��/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O Y/KOuO�O�O�/�/�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oQOcOmoo �o�o�O�o�o�o�o !3EWi{�� �������/� �o[oe�w������o�� я�����+�=�O� a�s���������͟ߟ ���'�9�S�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�K�9�g�yϋϥ��� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�C�U�_� q��9�Ϲ������� ��%�7�I�[�m�� �������������� !;�M�Wi{��� �����/ ASew���� ���//+/EO/ a/s/�/��/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? O#O=/GOYOkO}O�/ �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo5O'o Qocouo�O�O�o�o�o �o�o);M_ q������� ��-o?oI�[�m�� �o����Ǐُ���� !�3�E�W�i�{����� ��ß՟������7� A�S�e�w��������� ѯ�����+�=�O� a�s���������Ϳ߿ ���/�9�K�]�o� ���ϥϷ��������� �#�5�G�Y�k�}ߏ� �߳����������'� �C�U�g��w��� ��������	��-�?� Q�c�u����������� �����1�;M_ ������� %7I[m ������� )3/E/W/i/��/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�? �?�?�?O!/+O=OOO aO{/�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ O#o5oGoYosOeo�o �o�o�o�o�o�o 1CUgy��� ����o�-�?� Q�ko}o��������Ϗ ����)�;�M�_� q���������˟ݟ� 	��%�7�I�[�u�� ������ǯٯ���� !�3�E�W�i�{����� ��ÿտ�a���/� A�S�m�wωϛϭϿ� ��������+�=�O� a�s߅ߗߩ߻����� ����'�9�K�e�o� ������������� �#�5�G�Y�k�}��� ������������� 1C]�Sy��� ����	-? Qcu��������� �$ENE�TMODE 1I�^� +   (/�:+
 RROR_P�ROG %*%�}/�)X%TABL/E  +h�/��/�/�'X"SEV_�NUM &"  ��!!0X!_�AUTO_ENB�  D%#U$_N�O21 J+9!�2  *�u0�Ju0�u0�u0(0+t0p�?�?�?N4HIS3�
 G;_ALM �1K+ �u< +�?/OAOSO�eOwO�O�?_2T0  +s1:"�J
 �TCP_VER �!*!u/�O$E�XTLOG_RE�Q�6�E9 SSI�Z)_TSTKFY�c5�RTOL � 
Dz�2�{A T_BWD�@p�P<6�Q8W_DI�Q7 L^G48$x
?"�VSTEP�_��_
 �POP_DO�h_!FDR_GR�P 1M)B1d �	�Ofo: W`�������gl�pw�q�����I �����fWc�o�mW`C}��XB��FCd���A��BֿځB�;��mB�)��A��B�H�
A���A���m�o3�WB{f��p/�V!A.�>��Β� 
 Eǻ� �b�pr�wN�B��8�#�\���m`}dC��N���B�{���m@7UUT��UTF�Ϗ�j��s���m�OHc�EP]��O���#M��*�KA����m?�F��:6:N�r��9-�z��m���+����m���u(<!�����z�;�+FEAT?URE N^�P�>!Han�dlingToo�l � mpBo�Englis�h Dictio�nary�
P�R4D St�ڐard�  o�x, Analog I/O��  ct\b+�g�le Shift��  !*�uto� Softwar�e Update�  fd -c�m�atic Bac�kup�IF O���groun?d Editސ��g R6Ca�mera3�F7�P�art��nrRn�dIm���psh�i��ommon calib U����n����Moni�tor�CalM��tr�Reli�abL��RINT�Data Acquis�Z�Ϡ~C�iagnos���0�<�almC�oc�ument Vi�ewe�\���C�u�al Check Safety���  - B�Enh�anced Us抰Fr���8 R�5�xt. DI�O �fin� (��@ϲend��Er�r�Lm� D ph^���s	�EN��r.�հ �P�rd�sFCTN /Menu��v8����m�FTP InN'�facN�=�G���p Mask E�xc��gǱisp���HT^�Prox�y Sv��  V�LOAאigh-wSpe��Skiݤ/ ef.>�Hf�ٰ�mmunic��o{ns�
!
���urE�'�7�rt �F4�a�con�nect 2;�I�ncr`�stru����� SpK�AREL Cmd�. L��ua��O�AD*�=�Run-;TiưEnv� �yD;�(�el +��]s��S/W�.{��Licens�e����
����og�Book(Sys�tem)蔭�J�MACROs,~��/OffseS��Z�MHٰp��� j;73ΰMMR���l�35.f��ec_hStop��t��R� ize*�MiL��O� 2�7�x���0����miz��o}dM�witch�h���a�.�� v�ދ�Optm��49����fil��O�RD��0�g�� 8�496�ulti-�T������CPCM fun,�^�.sv�oO�Ğ�� �^�5�ReKgi��r��	�!2��ri��F�  H�59k�1�Num �Sel*�  74� H��İ Adjyu���adin���O� ,[���tat	ub��\У��������RDM Rob�ot��scovej� �d em(�:ٱn� SW��Servoٰs�����SNPX b���1��g P�Li�br���1ăڐ 9� ɰ.3�0g o��tE�ss�ag� f�"�@ e����"g���/I_�
�I�TM�ILIB���� P Firmn���^�F�Acc����0���TPTX���5w10.� eln����������H57�3�rquM�imgula��� 2�7Touz�PaxѩE1� T��6���&���ev.��IU�SB po����i�P�a�� 0\s�y nexcep�t��3 <� \h5�1 ����odu�V#��9��Q�VxN�k"6PCVL{&��^}$SP CS�UI�d���+XC���auҠWeb Pl���t? �#S ��\"	2�������S��&ު�V?8Gri=dplay��&�� ��8�-iRb".�� @ � R-20�00iC/165�¦ d+�+�lar�m Cause/�1 ed�<0:�As�cii����Loaqd��V4�3Upl�0�_CycL�c�m��ori����FRA�[�am�) tdt���NRTLi�3O}nݐe Helݨo 542*�PC`��4�`�]�1tr�ߵ48��ROS Ethv�t[����10\ҠiR}$2�D PkߵDER0>1�E����of�A��,ΰ�FIm��F�� �z��64MB D�RAMު�@:�9RF�ROA[�Cell03� ����shrQ
�B�Zc���ÍUk�p�� pide�Wty2L�s��|0\z�!C�tdѰ�.��@"Emai��li���+С\�� R0�qZ$GgigE�N�4OL�@Sup"��b�W3oa�~�cro�������4��QM��Fau�est�A>�j�� myiH9.dVirt��0W��0{&ImM�+T����}$Ko�l B�ui��n�յ'AP�L�&��MyV6� "\�0�*CGP�l��փ{RG�'p�{SB�UW�RQ�)K�&c�m\:��z��fX�)Oؒvõ(TA�&sp	oҠ-�B�&��
 I�f\E P�+�CB'f�g-��&" 5 �E��sv�b��Hvv�3��S_k��TO;�-�EH�f6.
�EN�vfx_z�)�V���tr>�)�hZ%.�F��& � ��r���*�G��&���њr����Hx��РJzCTIAc�pw4�LN�1�Mr�" #[��g�"��M�-�P2�~Tp�@����vxui�-�S�&�S�&�*4��W��2.pc�)V�GF��fxwʪV{P2AU \fx����N�if�u���"�in��VPB����)��s�D��*��a<s�F�5 M��s�I��c��{&Traİ��U~,p  ��<��2���RDp	�N���HY���p��-���H���Øp)����� �ϭ����yħ���rд��Ϟ�í4+���'�9L���ӎ��yy�9ӫ�c3ߞU��B�O�q�u���kߍӍSyy*�ߩ�\Yy�ߞ��k�W���ӄ��Yx����:�y	�������5�o�e/�Q���,�K�m��yg��^~��Ε�u�2��A��y������F������y�)���|�����1�m�.�<+�M��8G�i��7n��c���1�� ����W<�����7�{�����6�Z�������uk��[�|��!��?�ϔ��i�B\����_���{�x@.��wrst���B��� H68��@H�)T@J�EEND9I?��tql[}�
_�w�P�T�Q (��I) "���PA���T��/��85/A#b s;/�C/U/�,q�/�B�Gp�/�#��/�"3�6�5�R ?!2epai?5!:/Y4W���%INTo?e?_.�q�?4)��?�2pas2g�?�F O�?fA�ad6?��t Z�UD2gunOOqC5#33R?�D�0u�O�/��Mcm���OO�LNT�?��P_�Ĕ�0_0QR7�L_�Cfi._H?8_,_f'R50�_�S�AF-F�_�7�w.vo��_�_8�/�dM Cbo���o�bvrEo��paa��oaD�@�osF-A�S-sS�p'Is(8�PCesXPL�O�tslo_�ut\a�O�h%afvh%- B ��/����C�$��srp�?@_�?`w�"}�bA�����h�`���]T�ˏ�sgch��os�t��CG\s�;��us�?���Sg��/�G J����G�Dǟi$"�o�gdiʏ!�fd���?�h%J64S��Tut �o�O�?s����F�_夀���E�0���D`!��)�NO4E�O�i$II���iwjOl�ž0��>�?*�lb
��V��vjr/��
���7���ϥ�_�?zG7\ 2O�EG��Ϲ?���1՘ ޯ��_d�oi�8 ��c�50�>�x�Ͻ�"Lo�h%����dj9�﴿ƿؿ�c�� up9�C� j9�{�E��L��Ek, B串����oS_e_�&p/��O}�j94J���duZ��U��=d`;�����8���r7�Dhu���;]m T��������f�a���M���0�P�-4r V���O" #S�dwcL�P�in�`�a�?f& HTuRef�&��
�?hc�g�qr"��q.JG"�erM/��/ �/LsRA^��uH71�/��tCK�/<eTXP�/?i�k1/m5k.f���riR�eHG�/�/ cr�N'HGRf?L�iY�7�2hOuX��H\mO�� oρ�;H��DD@�O�� *�<�:I�?�?��d�R�η_ hd�ghg`OO�_���gmh�_h�m��XO�o|O�O�o��O\/�o0�f�gm �o`��`e۠;i�ov��yt��"��uRc60���#tmo�_�#1��fd r,op7��_�����lp>oh��冬'~ ߏ�dgts���&dޏ�/�o0�o
�J?<�vrF���cv.R���Ɵpld�56�%4�0/���greeK�m�XP)�fKCO*O|%56?��OZ� o~����E$i�o����jߠ���l ̂���OR��LOFvod��_IF��$��� ߪ�DߦX!B� Uc�e��t�4 ���(	M�O�5)e?Ƕ/���`1?Q�D�uk� '�|����`�boto�����-���6�p�eS ��on*���^� lB'����Տ_�q�_�rdk��4f��C( ҿȿ¯ԯ������̟p�����
I���571��t�ad�i39Tar��l�o�fk�������vPå@� PJ��|*���������e�t�4epg���ed��� E�5�RI�  H5�52� 747�2�1�pWelRK78�,� �0E�TXJ614���ATUP � wmfh 54�5�p�"6�pk��VCAM  7�\awCRI�@ ED" G UI�F)!28  j�CNREM�`��63�a�SCH�  4C DOsCV� CSUi��!0 D sEgIOCE�54�n#R694 we!!ESET=S#!3!�a� 73!fanu�MASK��OPRXY�_"7� ��0�OCO��"3�=P[�#"�ER J��" 7�!!J77�4#!39�  Eq8�G1�LCH 0#�OPLG%J50�00#MHCR)%P�S�17#MCS 4pD"�04 O#J55 �[#MDSWe!Y1M�D#1s#OP#1#MPR$07�0w"0�#8�  �#PCMX �#R0A�#� &�00��#� ( �&0�$50�( �#PRS� 3Js6903FRD@ �02RMCNy�n�dM�93 �SNBAA�80�0�@HLB  "�Lo�SM�A0 �(Ww"4 onitz#!2  II)��TC [#TMILpe �B�`0"K3�@�TPA� �QTXna�t\j�@EL�B&M250`0/D8��$�78�mon�19�5d SD95\FUEqC 0OP� UFR@ ���;!C@ \�@;!O:�0pt"VIP�@#� I�@0�!CSX�� �#WEB �#H�TT \stB2�4 �#CG�Q#IGޫQtopm�PPG�S!��PRC�@SH�7���w!6( �8���![�R RBB- sCi�B01rogw!f#IF#"098-!�!` �@�A64�(AaNVD�!Ld�1h 6a68( c�`d S{R7c!te.p� �0kaч@�bc`� CCLI$0?�sb$c9G �MS�"5a�` - �A� STY�@al� �@CTO �CJ�NN0J98�O�RS�0G��b�g �J�`OL�1Abn�: SENDu�to��!L�Q���@*r#S�LM� 8�"FVRn� MCHN0CSW!�SPBVP�� P%L� ds �qV$0�c�CCG $p�aCR҄0
Np�QB� 87�.f�QK� j70�*`�p�0'3CSqToo�CTQ���q�TB�P�N��@n$;pqC�@�Q#�� �p,#�p ��. %�$0h7#%� `8D#TC� QSQ"TE� [#m�, �tTE� gt"m�P�TTF�Q[����@�#CTG�Q�"���@ί#CTH `�TTI�@#CT'Qeqs�PCTM�@SC�$0xgS��0bodyq=P�@  ��� O�1� d��q�aus�a9��P[��qW `@06; GF� `8�V@VP2@ 6#23R i��@j?�g�R `n�g�B `" �g�D `��g�FX m;na"PVPI��+ �G V�!#V	`  23�RVK�@Np�@�CV�Q31�93{4.�vo R�erne땗�����i��r���h����A���37� ��"�\srv�����b�3b�- Sr�B"0���A�J935땿B�/5 (S�O���g �1�1�R|��j93땷b��ENz�5�� awm�{SK� Lib� �������� ���	 �"|�h�h��#��b�wmsk"�nE����q����pyE�  ���!x�02�t Fuï�բ6ۯm��uji%-�I&���8k�� 8!�Ń�땼P��2�p2�2�Mai'�on��_�/r�;pڦh;�;�G��_r���!v��4\ֶORC�ֺ+�5�� "T¦T�P��hQ�652�10��4���<�xk������ߦ�t�P��QrxֶSB�� ch_�����)�t!0�B�"̿ h�h땇�;���c��� ���������>�Rp� \toֶ3���#cl�W��2p�"� ���������F� ���b� Qt�a�϶0�t��ܐFsȒ�76t�p�t	� Ad����582��ob�|g*{�\a���FMQ ���A�mi1gֶ�I�or�w�I�j�rfm��F�c���@1�EYE&~� w���R����4�K2Х70.�E�ld,�C�� 1PTP]���..�"AD.�F�&83 k���ask���"�`4���۳dֶےv��ER~�7 R�ƀ�/�T�?)�e�rv�G?Y?k?}?�?�?ӹapa��	d��h��r�4�M��te��"��79!J�d/���G�p�ac�T��<�6�b�/� QO��$v�c>�,@Vg����e�YW��5/� BJ�h���R5:�d��Ɓ0�@��I_�raaj��e��he}ǔ$`��5(Xa�@��eqt榻�1Otdj��h,�_h�\	UI�/k�jo�FO��`^���aF��r��qW65q���K �'6ڦus W'�b,'��'?��n��MFR��;]�blf�ǯ�fr>���w�p�/�,��_U[ǀ�мn�x'_i� {�����O���pJ���X[@�o�in7L��O�9�\^ �� R����+mi�2״h �j��҇- �f�nt >�MA� H�I  �H5529� (�Cߑ21��le�R78�c�ߒ0�AcaJ61�4���0ATUqP�����545�t�-fl�6yE=�V�CAM�tFLX�CRId���o�U�IFULX �2u8��mo�NREu'���63��WQ��SC�H��Cn�DOCV��gϠCSU1�cx�r�0$�;EwIOC%tx\c��#54�oQ��9T�;��ESET�Temo�?�S�/��7S�{�M�ASK��70��PGRXY�T�`��7�ú`�OߐOCOe�\B?�3�ô`>��0{��?��|�-��on G?�39!'ߑõ� H82LC�Hd��@IOP�LG�tCGM?�0x��GЎ�MHCR�Gbo�S�/1_�CS4�7cgm��50T���?�5$�[���MDS�WMf.�D�����O�P��X/2L_�PR��K�����{����883n�CM��0iA,��0�Ő`~�=5#�\h88��+�?�D���.?���4J��0D�3��o�S4�����9��,i�FRDd�/2E/���MCN5�H93��K�SNBA�U"�R��HLB��SM�՛ñ�T���J52��SaߐTC4�\�T?TMILe��Pt���A|�TPA�^��TPTX��5��'TEL�ԫ�0䴈P���8�˳���K�9�5����95��88�8��UECd�rt �UFRd�__��Cd�2e-�VCO4��VIP�;���I�TAX~�CSX8�����WEB4�����HTT4�ka��2^T�2M/So�G#��QIG��< .��IPGS=t\rxFO�RC��aߐ7��/a��6D�s@>�R7 #��!��Oq�Ҥ��P ��Ҷ;�A���KÑ�$��0 "��4����N�VD4���#�Adaep��8D���68��ƻ�R7���P��D0���a��o�bܠ. CLI��l\-C����CMS�'��4�d; "ްSTY�[�CTOT�tl��N9N����ORS4�;��1 ��ltiΰOLS�( E���0�T���EL��6�@���9@ ���LM4�HV fo�VR���CS��wshc>�PBV4�쫁/�PL�
APVust>�CCG�4��0nCR�4 �H5��B���K�H573���?�<���\cms�#�7st.~TB���(! ��7�C�ԓ�<?"�awsh?"���I0?"��3�TCpd�K�A 4�\sl"AEĤpP��� 4�C[��"Ԥ8c��"4�(��CTF��c��"�n��CTG�73m#YG�THd�h� ��I��K�CTC�5�9m�CTM�5M𔴻�Q0��re\g�P���12��0�4�����%S��1]3MCTWd�9[@�_�GFd�SE]�P2d�t+��2�ա �2nd�ell��PBd�I���1Dd��a�1Ftap VPILd���CV�!Vq�:�UA��CVK�ۣ�CV#�core L���H"�Hp!�HK"�Hatc�J�H��4�I� �IL0H �I�2�H��H+2�IL��Y4=�H���Ie\1a�I�2 Z93�I{ �H�@NZ+��H 1��K#48�Z<A�Ht{�I l �Z;"�O�Fs\!�H�k"�H{"@o�F[�PZo�Z���J��Tok�РH��H\��Il�Z���Z2=[ng-[gT�oo�I�p�j(�njr�obt_�Xbt.�JL� iur�o�I� �i�!��F��POz�ling�j��y���Y"r^zۢ�I�p��Geat^j�]��Z��_je�����_��lkҠHm,��H|��Z���A�I  �_�s  ���Gvhm�J�{�svnj���H49�\�J�@L�Ij74u9{P�Zt\jNj��@_"g.pjmc3al�0�fu�J��^zhm-��_bg���o��\ͫ �1�H! �j��;����MT "�(Cu�zk��bg�ft�JlpX���GgCT"���Gfc]��˝26\fߟ�9C26�l\� Ίup�>m��;�Mul?��Q��7\^�K���7`-[˝���_�61Nj748.� H- �H��@R_�L^ziPe0��K�Я�F8\}�}�`����Ћ� � Rk,�ticMoj+@Oo�Qxs-@�"�3�CS� j+}LB-[5 9HNj+� co~�L�d�z��f�k˝lb��jll����-˜�k�/�.���LЎ�kipJ/�on,�J\A��]8�SK"�� ��wuto�o B��X����kwm� �o��Htp�ʜ n}��#ex-�˝��x���%a^jlL�je�식	i��a��/���{rej�1�o,�Vor�zR�����e T�Z[��[lc�lN��߭�SOžG3ZD��to�{+BΠH643N�`�SG/o��sg�a�Utui��;`�J��`��;�ndm�ndi N�{/�/�/�/�/�/�/��/??/?A?�?��r�iΪ! -Kj95�0/�n �zk]8915n/�O�t �Z���wsg�K,�>��i;ag� SGJ����ogu���KO]Lstw>_@	J64�:1�s�{F O>ګ#cdݛ��`3_��Yr-��N74�y-��3��RINnzlly��(m^���L����sgc�zI" #p?
+�oߡ\tw/� ��0.�@�"���f�_ʯ[y�Kmm�K}dc�t^�t]�+�
PR�ZWCHK
k, �;;`y<p��lK����LN*R85j ̛@_jR ���ti�N�g WJhecdN�L�F����wlZw|*�dat��Λ�greN��o�  STD��r7LAN-G�Aoc�e�`���Q�7��R87�0�{��8 (P�ogge����!�58\�PAcTTs�� �t\�N�c "B�@V�<�1�patd���O���������{q�
��5�a�p[�m�\q㕻�7�\aw��@�a��p6�����<ϯ�gmon���d��0�B�m�;A���\ ö��K�I�MH{CR�51 H��B��g\o��@��R]Ǐ H54ۿm�<@E����;!�����om�m�;a��R�|�N㕬0F�C��W�P�)Ai6�� Fƫ�{��itx�#{ ��icaio����De6��eve����72 �R�@RƜPg��ad�l��nt��K�RBT�tOP�TN`772'�CTK"'�g�(䔠�)� "AZ'�;q'圻q'�tzn&�{ E�'�Ama��- M�u��ncInDPN�������O872��|�d��(��������#����masy��y "�M��o��䃲��et����\p1�����\ 2��f���lZ����lp���9���`��+ V��ail��?������䓢��zd�<�k`���73.f��ir�dg��- i��ep\ ����� S0j�021"�1W ��(��`�4�� (i��e,"� "���+���/core_�I��l`aF��AY��AB���@����H�����AB;IC��Par;�M�ai������<� ;c\�ITX>����  ����1���g Jclib��ShiW�4��� t994\�V�SSF��� tt\{j9�f "O�pw� t��$%ini�/��pٰ t�5G�&�,� t\vsR&x�Lx�%w� tamclS/+ref.�%#� t	j��%m�� t[A�&�4\z�/�,z_v��%A�%�a�%_ol�6��l% �%end��/<c?.?@?R5o�[?m>�6�/�dshf�/+trt�?<O<AE�'F  !�G��$%��5vi�6���6� J92�F3��%2'5 (�%�@e&�Px�%k�4O dnwzFb��T�&`�XEpn�&|g��? nw\n�?&�,nd�V��N;XnF� j���%se�V I/
&�q&фU�n�5r w�%/F� X�F�_�rclR&0\p,w/Y�90�Eo`/:"5Of "U//A+dprm�%g¨%�XCrsu/kmS�T_ L`�6/OŔpM�LO�j��`nO1|h�ODnon8�|YCwrpR/�lp���E<�Pe\ga��Krgas�o�k�b�f�v��4xtfL�?m$ra�o�la00�omk�_�TamN6+�p4�`'9K0.v�W�ې�%�@�Ft��XE �sV��ДJ737�%|*�%,P���hB "+��Kwcf�F& I����998�vtomzFut  vV�_	o;�YC���:#8\F&�Y/� 0��f��deb^V��$@�0zFؠ"��g����<9\�&��9�Wrl}  �su"�st�G`��X �f� U (�fagn�F PzFϜ�V�ia�TX����v�d��w��g��HzF- O�W CH� �$G723�F���E(Aπÿտ2蚽Wc��Ws�vF& S�W�JR64��_�RVo RV���ӊ��vt�M\�etF�XoN�o�Fr ��x���+�1T�F?zteR� J58�O�  34	Wglea,�%,�j�Dq\t"���zFwIta1lUT�A�VϜ�gw韗Ma�d�W�Oa���6d �M��e�FT��90� H�%NT��R6�9������ir\�ʆMIR��ӊen�ʆv���F|�3��ITCP��Ta0�p����(MM7G�eT�o �\tpʆI��YBbusJ׈�m��I�@zFȀ��F�����/:��W�'g, ��4`�R_(!sw�&s_YC6c7\JF��Tf_�����Dfw��W��4a3chg��a96_���� _���_rV�% 99YA��e��$FE�AT_ADD ?_	�����?  	�$YA //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o #5GYk}� �������� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿�������DEMO �N�   ��*� �2�_�V�h� �������������� %��.�[�R�d����� ������������! *WN`���� ����&S J\������ ��//"/O/F/X/ �/|/�/�/�/�/�/�/ ???K?B?T?�?x? �?�?�?�?�?�?OO OGO>OPO}OtO�O�O �O�O�O�O___C_ :_L_y_p_�_�_�_�_ �_�_	o oo?o6oHo uolo~o�o�o�o�o�o �o;2Dqh z������� 
�7�.�@�m�d�v��� ����ƏЏ����3� *�<�i�`�r������� ̟����/�&�8� e�\�n���������ȯ �����+�"�4�a�X� j���������Ŀ�� ��'��0�]�T�fϓ� �Ϝ϶���������#� �,�Y�P�bߏ߆ߘ� �߼���������(� U�L�^������ ��������$�Q�H� Z���~����������� �� MDV� z������ 
I@Rv� �����/// E/</N/{/r/�/�/�/ �/�/�/???A?8? J?w?n?�?�?�?�?�? �?O�?O=O4OFOsO jO|O�O�O�O�O�O_ �O_9_0_B_o_f_x_ �_�_�_�_�_�_�_o 5o,o>okoboto�o�o �o�o�o�o�o1( :g^p���� ��� �-�$�6�c� Z�l���������Ə� ���)� �2�_�V�h� ������������ %��.�[�R�d�~��� ����������!�� *�W�N�`�z������� ���޿���&�S� J�\�vπϭϤ϶��� ������"�O�F�X� r�|ߩߠ߲������� ���K�B�T�n�x� ������������ �G�>�P�j�t����� ��������C :Lfp���� ��	 ?6H bl������ /�/;/2/D/^/h/ �/�/�/�/�/�/?�/ 
?7?.?@?Z?d?�?�? �?�?�?�?�?�?O3O *O<OVO`O�O�O�O�O �O�O�O�O_/_&_8_ R_\_�_�_�_�_�_�_ �_�_�_+o"o4oNoXo �o|o�o�o�o�o�o�o �o'0JT�x �������#� �,�F�P�}�t����� ����������(� B�L�y�p��������� �ܟ���$�>�H� u�l�~��������د ��� �:�D�q�h� z�������ݿԿ�� 
��6�@�m�d�vϣ� �Ϭ���������� 2�<�i�`�rߟߖߨ� ���������.�8� e�\�n�������� ������*�4�a�X� j������������� ��&0]Tf� ������� ",YPb��� �����//(/ U/L/^/�/�/�/�/�/ �/�/�/ ??$?Q?H? Z?�?~?�?�?�?�?�? �?�?O OMODOVO�O zO�O�O�O�O�O�O�O __I_@_R__v_�_��_�_�_�_�_m  h$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ ����"�4�F�X�j� |�������Ŀֿ��� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�t߆ߘߪ� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: L^p����� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲���������>�  �� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZl~���� ���/ /2/D/V/ h/z/�/�/�/�/�/�/ �/
??.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo Xojo|o�o�o�o�o�o �o�o0BTf x������� ��,�>�P�b�t��� ������Ώ����� (�:�L�^�p������� ��ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ�������� �*�<�N�`�r߄ߖ߀�ߺ����������	�,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oi��$FEAT_D�EMOIN  Vd�D`�`,d_INDEX9kHa��,`ILECOM�P O����zaGb'ep`S�ETUP2 P�ze�b�  �N �amc_AP2�BCK 1Qzi  �)h�o�k%�o`}`A e�om�o� �� V�z�!��E�� i�{�
���.�ÏՏd� �������*�S��w� �����<�џ`���� ��+���O�a�🅯� ��8���߯n����'� 9�ȯ]�쯁���"��� F�ۿ�|�Ϡ�5�Ŀ B�k�����ϳ���T� ��x��߮�C���g� y�ߝ�,���P����� ����?�Q���u�� ���:���^������ )���M���Z������ 6�����l���%7 ��[��� �D@�h��i�`P�o� 2�`*.V1R`� *c�`����JPC�|�� FR6:�".�4/�TX`X/ j/�U/�,;`%/�/��*.FM�/�	���/<�/<?�+STMG?q?��]?�=+?�?�+H�?�?�7��?�?�?EO�*GIF OOyO�5eO"O4O�O�*JPG�O�O�5�O�O�OM_�JSW_�_� �Sn_+_%
Ja�vaScript�_�OCS�_o�6�_��_ %Casc�ading St�yle Shee�ts0o� 
ARGNAME.DT_o
��0\so1o�Q�d��o`o�`DISP*�o�o�0�o7�e)q�8�o
TPEIN�S.XMLg:�\{9�aCust�om Toolb�ar��iPASS�WORD.�F�RS:\�� %�Passwor�d Config @����������� r�����=�̏a�s� ���&���J�\�񟀟 ����K�ڟo����� ��4�ɯX������#� ��G�֯�}����0� ��׿f������1��� U��yϋ�ϯ�>��� b�t�	ߘ�-߼�&�c� �χ�߽߫�L���p� ���;���_��� � ��$��H����~�� ��7�I���m������ 2���V���z���!�� E��>{
�.� �d��/�S �w�<�` �/�+/�O/a/� �//�/�/J/�/n/? �/�/9?�/]?�/V?�? "?�?F?�?�?|?O�? 5OGO�?kO�?�OO0O �OTO�OxO�O_�OC_ �Og_y__�_,_�_�_ b_�_�_o�_�_Qo�_ uoono�o:o�o^o�o �o)�oM_�o� �6H�l�� �7��[����� � ��D�ُ�z����3� ԏi��������ß R��v�����A�П e�w����*���N�`����֦�$FILE�_DGBCK 1�Q������ ( ��)
SUMMAR�Y.DG����M�D:3�s���D�iag Summ�aryt���
CONSLOGi�L�^��������Console log�����	TPACCN��R�%:�wς�T�P Accoun�tinρ�FR�6:IPKDMPO.ZIP�ϯ�
����σ���Excep�tion ߱�_�MEMCHECKm��Կb����Mem�ory Data|��֦LN�)n�RIPE�\�n����%�� Pa?cket LϺ���$SA���STA�T�����ߋ� �%�Statuys��<�	FTP�����r�����mment TBD���� =�)ETHERNEU���B��S�����Ethe�rn(��figu�ra߇���DCSVRF���������� verif�y all٣M�(��DIFF�����/di�ff�PB���CH�GD1�x�c �FQ&��	�2�� 85�YGD3���'/ �N/��UPDATES�.m S/��FRS�:\k/�-��Up�dates Li�st�/��PSRB?WLD.CM�/����"�/�/�PS_ROBOWEL1���:GIG�ߊ?/��?��GigE ~��nostic*�~ܢN�>�)�1HADOW�?�?�?�5O��Shado�w Change���٤&8+�2NOTI��O"O�O���Notificx��\O٥O�A�� _��2_կ?_h_���_ _�_�_Q_�_u_
oo �_@o�_dovoo�o)o �oMo�o�o�o�o< N�or��7� [���&��J�� W������3�ȏڏi� ����"�4�ÏX��|� �����A�֟e��� ��0���T�f������ ����O��s����� >�ͯb��o���'��� K��򿁿ϥ�:�L� ۿp����Ϧ�5���Y� ��}���$߳�H���l� ~�ߢ�1�����g��� �� �2���V���z�	� ���?���c���
��� .���R�d�����������$FILE_�� PR� �����������MDONLY �1Q���� 
� �)�@_VD�AEXTP.ZZ�Z��p�G�L6%�NO Back? file !��U3�M��7� ���G�&�J\ ����E�i �/�4/�X/�e/ �//�/A/�/�/w/? �/0?B?�/f?�/�?�? +?�?O?�?s?�?O�? >O�?bOtOO�O'O�O��O]O�O�O_(_��VISBCK����*.VD)_s_�@�FR:\BPION\DATA\^_�R�@Vision VDt�_�O �_�__o_Ao�_Ro woo�o*o�o�o`o�o �o�o�oO�os� @�8�\��� '��K�]������� 4�F�ۏj����̏5� ďY��j������B� ן�x����1���ҟ�g���MR2_GR�P 1R����C4  B�O�	� 
������E�ˀ ֯�r���OH�cEP]��O���#M��
�KA���?�&�r����:6:N=�R�9-�Z���A�  v���BH���C`}dC��=N��B�{��r����пὫ�@UUT��U����/Ϫ��>��>c���>rа=ȫ��>i�=����>����:���:��:/�:6)�:��~ ϗ�2ϔ��ϸ�������z�_CFG =S��T  �a��s߅�0[NO ^��
F0�� ���/\RM_CHKT_YP  ���O�h���������OM���_MIN��L�������X��SSuB7�T�� ��5�L�,�U�g����TP_DEF_O�W��L�����IR�COM�Ѝ��$G�ENOVRD_D�O��	��THR��� d��d��_E�NB�� ��RA�VC��U�UQ ��Υm�X��|��������� � �O�U��[��O�x���⾥8�:����
,.  C�x �h�������B�ϡ�����n�.!�SMT'�\.����+�w�$HOST�C7�1]K[̹Y��� MCL��MI�  �27.0�1�  e}��� / *�1/C/U/g/�!/�#	anonymous�/�/�/�/�/"? L��8;{ }/j?��?�?�?�?�? /�?OO0OS?�?�/ xO�O�O�O�O?UO+? =?_QOs?1_b_t_�_ �_�?�_�_�_�_o'_ ]OoOLo^opo�o�o�O �O�O_o G_$6 HZl�_���� ��o1o� �2�D�V� h��o�o�o���ԏ ��
��.�uR�d�v� ������?������ �*�q����������� ݏ��̯ޯ��I�&� 8�J�\�n���ǟٟ�� ȿڿ���E�W�i�F� }�jϱ��Ϡϲ��ϋ� ������0�S�Tߛ� xߊߜ߮�����+� =�?��s�P�b�t�� ���ϼ��������'� ]�o�L�^�p�����~/ENT 1^��� P!���  ������*�� Nr5~Y�� ����8�\ 1�U�y�� ���4/�X//|/ ?/�/c/�/�/�/�/�/ ?�/B??N?)?w?�? _?�?�?�?�?O�?,O �?ObO%O�OIO�OmJQUICC0�O�O�O_�D1_�O�O�V_�D2W_3_E_�_!ROUTER�_��_�_�_!PCJ�OG�_�_!1�92.168.0�.10�O�CCAMgPRTGo#o!7e11@`noUfRT�_ro��o�o��NAME �!��!ROB�O`o�oS_CFG� 1]�� ��Auto-started��/FTP��~q� ��F������ ��9�K�]�o����&� ��ɏۏ�����Wi {X����o�����ğ ֟������0�B�e� �x���������ү�� �����Q�>���b�t� ������q�ο��� �9���L�^�pςϔ� ��������%��Y� 6�H�Z�l�3ϐߢߴ� ������}��� �2�D� V�h������������ ���
��.�@��d� v���������Q����� *<���� ���������� �8J\n��% �����EWi {}O/��/�/�/�/ �/��/??0?B?e/ �/x?�?�?�?�?�?/ +/=/�?Q?>O�/bOtO �O�O�Oq?�O�O�O_ 'O(_�OL_^_p_�_�_�(�`_ERR �_z�_�VPDUS_IZ  9P^S@���T>�UWRD� ?EuA� � guest3V$o6oHoZolo~o��dSCD_GRO�UP 3`E| �Iq?YM �nC;ON�nTAS�nL�n�nAXP�n_E�o�9P�n�RTTP_AUTH 1a�[� <!iPendan�g�~@}9P�J�!KARE�L:*���}K�C����pVI�SION SET�`E��I�!\�J�t� �s����������Ώ���-���dtCTRL� b�]~�9Q
�`�FFF9�E39�DFRS�:DEFAULT���FANUC� Web Server����bvod L��'�9�K�]�o��T�WR_�`FIG �c�e�R����QIDL_CP�U_PC9QB��@� BHǥM�INҬ�a�GNR_IO�Q�R9P�Xɠ�NPT_SIM_�DO�!�STA�L_SCRN� ��y�+�TPMOD�NTOLY�!���R�TY8��&�9�hpE�NBY��cƣOL_NK 1d�[�` �����1�C�U�Ͳ_MASTE����&�OSLAVE �e�_˴jqO_C3FGsϦ�UOD���>��CYCLE�Ϧ����_ASG 1f���Q
 W�9�K� ]�o߁ߓߥ߷�����������#�_��NU�M�S�b�U
��IP�CH��j�O_RTRY_CN��Z<��U�_UPD�S����U ������g��θ`��`ɠP_M�EMBERS 2Yh��` $�e��>��HyɠSDT�_ISOLC  ����r�\J23�_DS��q���O�BPROC��%�J�OG�d1i���89Pd8�?�.���.�?�?�?OQNs��V����3W~������������POSRE���$�KANJI_�m�K�i�pMONG j�k~�9Ry� ���//�^�r��	k����9%Th��p�_L�I�l�kEY�LOGGIN���`����U�$L�ANGUAGE Y����� �!��QLG��lq�9R���9Px�p�  j��砬9P'03X��k���MC:�\RSCH\00�\��� N_DISP m��DAM�K�SLOCw�آD�z ��A�#OGB?OOK n����9P~��1�1�0X �9O%O7OIO[OmN�M0ɱ���I��	�5I�b�5�O�O�5�2_BUFF 1oؽ�O2A5!_�2�� =_?7Y_k_�_�_�_�_ �_�_o�_o:o1oCo Uogo�o�o�o�oe4��DCS q�= =��͏L�O-�1�CUg���bIO ;1r� ��s20������ ��1�A�S�e�y��� ������я���	���+�=�Q�|uE�TMl�d����Ο��� ��(�:�L�^�p��� ������ʯܯ� ����7�SEV��u=.{�TYPl���z�0����!�PRS���/|S��FL 1s�}����$�6�H�0Z�l�~ϯ�TP� l��i��=NGNAMp��A5�"e4UPSm0�GI��\!����_�LOAD��G �%u:%PLAC�i�2�3�MAXUALRMI�c�W�T���'_PR����3�R�Cp0t�9�M����3Eݗ���P 2u��� �1V	i�00���߭� 1��.�g�xU��� �����������8� J�-�n�Y���u����� ������"F1 jM_����� ��	B%7x c������� /�/P/;/t/_/�/ �/�/�/�/�/�/�/(? ?L?7?p?�?e?�?�? �?�?�? O�?$OOHO�ZO=O~OiO�OK�D_LDXDISA�����zsMEMO_A�P��E ?��
 b��I�O_"_�4_F_X_j_|_R�IS�C 1v�� � �O�_ ���_�_�Oo�o@o�_C_MST�R w:�_eSC/D 1x�M�4o�o 0o�o�o�o�o P;t_���� �����:�%�^� I���m������܏Ǐ  ��$��4�Z�E�~� i�����Ɵ���՟�  ��D�/�h�S���w� ��¯���ѯ
���.� �R�=�O���s����� п����߿�*��Nπ9�r�]ϖρϺ�PoMKCFG ynm�����LTARM_*��z�����и����6�>�s�METP�U�ӫІ�viND>��ADCOLXի��c�CMNTy� l�g` {nn��-��&�����l�POSC�F����PRPMl����STw�1|�[� 4@�P<#�
g��g�w��c�� ������������ G�)�;�}�_�q�����������l�SING_CHK  |߿$MODAQ�}��σW��#DEV �	�Z	MC:>WHSIZE�M�P��#TASK �%�Z%$1234?56789 ���!TRIG 1~
�]l�U%�\!�S
0K.�S�YP�6�9"EM_IN�F 1�� `)AT?&FV0E0X��)�E0V1&�A3&B1&D2�&S0&C1S0}=�)ATZ�#/
$H'/O/�Cw/(A/�/b/�/�/�/? �&?���/ �?3/�?�/�?�?�/�? �?"O4OOXO??�O A?S?e?�O�?�?_CO 0_�O�?f_!_�_q_�_ �_sO�_�O�O�O�O>o �Obo�_so�oK_�owo �o�o�o�_�_L�_ o#o��Yo�� ��o$��H�/�l�~� 1��Ugy����  �2�i�V�	�z�5���𰟗�ԟPNITO�R��G ?k  � 	EXEC�1���2�3�4��5�� �7�8
�9�������� ��(���4���@���L� ��X���d���p���|����2��2��2��2���2��2Ũ2Ѩ2�ݨ2�2��3��3�3(�#R_GRP_SV 1��� (��@@w��Y�=�N�4"⸿���1���R�_Ds�����PL_NAME� !���!�Default� Persona�lity (from FD) ���RR2�� 1�L6(L?����	l d��nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ�������B2]��� *�<�N�`�r����<���������� ,�>�P�b�t�����B�J  ��\  �  ���  ��  A_�  B��T�� 
��������  ������B���p���  C�H CH P E�z  E�� E_�` E�;%��Z�*�~ �  E��Fl�@&��T Ai� dx �H�x�	$Hx(d�dڭ�}` (d��8(x x$$y XHtd D (DD dpWwX��	X �vXHX���)/y�y (� !a��  7%E	��Em�Xw$%X8H$%P�� �/�/ �/�/�/�/??+?=?8O?a?s=F�r?�?�?�?�6��E���EA���2�����  ���?Kزd�3�4,O:IO\OjG��0��|MTCҷ'4� � W%��O�O�N  h�H�O�JA  A��C����_�OC_9W�  � TB�LY��
��_�\�@Q�Y=²CÈ�V�`HR0� ʒ�P( @7%?���a�Q?ذaر@��6�&س��2n;��	lb	 � ����pX��U�M`��X � � ��, �rb��K��l,K���K���2KI+�KG0�K �U�L�2o�E	O�n��6�@ t�@�X@I��b`�o��C�N����
���}v��#���` q�m�|�kQ?�
=ô��  �Hq�o`!b���9�  ��a� �B ���ذa�s�G��}2�m��o�q��v�O���E	'� �� 0�I� ��  � Q�J:��ÈT�È=��9�l��b@|��� }~�Q����RSD����N8���  '����p?��P�b!p�b){�B���?�CIpB  X���ذ��C�A�av/ � {��	�o�Q�IB P��8�����P��ԕرD �O���O���A�,�>�Š
�`l�1�	 �٠p��� p` rl`:GT  �t�?�ff{O��įV� �P����aa�,!�/�?Y)R�a4�	(ذ]�Pf����a\c�\dƃ?333-d����;�x5;���0;�i;�d�u;�t�<!� +}�oݯ��b�Sb��P?fff?��?�&��T@��A�#$�@�o[ ,ž�x�	�&f6�ed� g���Hd㯸ϣ��� �� ���$��H�Z�E�~߾�&eF��mߺ� i���U���y���2���E�0����y�d� ������������ �?�*�܏r�8�.o�� �����T�); ڿPb������0��P��A��T C�=�ϵ��Y}��2��������C��W�C�>= �` Ca���B����(!�`�<����bC@_;C�9�BA��Q�>V{�������Y���uü��
/��S��Q��hQ��A�B=ן
?h�Ä/iP���W��È�K�B/
=�࿣��Ɗ=�K��=�J6XK��r#H�Y
H}��A�1��L�jL�K���H:���HK��/0	b�L �2J���8H��H+UZBu�a?�/ ^?�?�?�?�?�?�?O �?O9O$O]OHO�OlO �O�O�O�O�O�O�O#_ _G_2_k_V_{_�_�_ �_�_�_�_o�_1oo .ogoRo�ovo�o�o�o �o�o	�o-Q< u`������ ���;�&�K�q�\������Gϭ���� �C�aɏ Ĉ���CVF������+b� ��Kc�f�� 
E�����T�ٟt�(t��g_�h۟��������N��������3lC�(�:�H����T�f��t�.�3��}����k����q'�3�JJ�����گ���4��"�]P̲Pf��� ����⟛�ſ���Ի�����/��?�{x?�N�u�  fUh� *ϳϞ������Ϣ�t�0.��R�@��X�bߘ�߆ߨ�)Z�ߺ� ? ( 5�	�߀����B�0�f�t�  2 E%p"�E[@��N�"BXC��%@ߏ��%������)�;��������������%n�n�%"T�%��Xc
 ��!3EW i{��������b*[��P�I��v�$MSK�CFMAP  ���� �^�����pDONR�EL  X��[��DEXCFE�NB�
Y�F�NC��JOGO/VLIM�d��]dDKEY��=%_PAN�"\"DRUN�+SFSPDTYw�x���SIGN�>�T1MOT���D_CE_GRoP 1���[\���/��?&?��? Q??u?,?j?�?b?�? �?�?O�?)O;O�?_O O�O�OLO�OpO�O�O �O_%__I_ _m__�f_�_O�DQZ_E�DIT�$UTC�OM_CFG 1��Q�_o"o
��Q_ARC_��X��T_MN_M�OD���$�U?AP_CPLFo��NOCHECK {?Q W� ���o�o�o�o' 9K]o������vNO_WAI�T_L�'�W� NT��Q�Q���_7ERR�!2�Q��� �_t�������A*��Ώ�d``OI�}�P�x :_�t��C+���XG���k)�70�������8�?��4�ӏ��|d�B�PARAMJ��Q����_�����s�� =��345678901�� � ���?�Q�-�]������u���ϯ����������7�ODR�DSPEc�&�OF�FSET_CAR8�PKom�DISz�K��PEN_FILE����!$a�V<`OPT?ION_IO
/!�аM_PRG %Q%$*	�ά�WORK ��'=� ��K�7"U�h��f�(�f��	 ���f�7����M�RG_DSBOL  Q������L�RIENTT5O* ��C���Z���M�UT_SIM�_DطX+M�V~Q�LCT �%���R_�$aQ�'�_PEqXh`��b�RAThg� d�b�r�UP� �5� � �`���߼�����$���2�#�L6(L�?��	l d'�O�a�s���� ����������'�9� K�]�o���������H�2>�����/A Sew�N�<��� ����1CPUgyH���P��� �  ��  �U�A� g B��PB�����H��  ����U�B�pҶ�����N�P �Ez  E�� E�` E���;(����Z��/���  E���''���@#�U��T�AJ(�� E!Y!a!)!m!Y!u)%�)!Y!E!�%E!ڎ$� ^$A!�	!E!a!�%%�	-Y!Y%�-58� Z 99U%E!�D!	$D%%E!Q481X291�% �)95�/W#95)%91m5�a!�5/Z7��Z (��8�1�<a1 EE	�(�Em�494X6�E9=)%E15��  |O�O�O�O�O�O�O�O�__0_B_T]FЀS_y_�_�_�Vh��� ��_�[��͔on��_=oKg�]�]&�'�4 � W1%po�oX� g��g��o�jA�A��c������o�o$w�
��tB�(~ΐ��r�|�` q�y�$��O��1�'k�o'��3�`���0��P( @ED�D��q?Q�C�Z7}��o�  ;�	lD�	�u� ���pX�[�2���X � �? �, �W�ΐ�H��9H��H��H`��H^yH�R��l���_����	�#�B#�B C4ӄ����c�9���
=���� �������cBz���{�a�m�� �b�s�� �q���g�2��챏Ǒ�ٖ�o����e	'� �� �I� ��  �q<�=����9�K�E�@�a�g�b����������E������N�� C '۰��Ɓ"�B�@Ղ��т6��� �?  ��C�a��!	ŀ~��p=�Bp���Н����px����D ��o޿�o��&��6#�5�Ю`Q��	 ٠U�*f� U� Q�:����#����?�ff0\o�ϩ�;� �p�����F�8� ��?Y�
r��q=�(� B�P�K�fɆ�A�A���?3�33��Ł;�x�5;��0;�i�;�du;�t�<!��y�������t���r�p?ff�f?x�?&���@��A#	�@�o[�	]��� ���uI��wh���-� �ϝ���������	� ��-�?�*�c�u�L��� ����4�V�X����EjPf��^I �m����  �$��W��� ����9��/ / ��5/G/�z/e/�/�/0�/�/�`�A��$�t�/ C�/"?�(d��>�?��Pn?�/�?�}?��(��W�?C=�@�` CT��?đj4�j0i1A@I��!���bC@�_;C9�B�A�Q�>�V`.È�����Y�uü���
�?�3��Q���hQ�A��B=�
?h���iOJp��W���ÈK�B/
�=����Ɗ�=�=K�=�J6�XK�r#H��Y
H}��A��1�=L�jL�K���H:��HK��O��@	bL �2�J��8H���H+UZBu �?F_�OC_|_g_�_�_ �_�_�_�_�_o	oBo -ofoQo�ouo�o�o�o �o�o�o,P; `�q����� ����L�7�p�[� �������ȏ�ُ� ��6�!�Z�E�~�i�{� ����؟ß��� ���0�V�A�z�e�Gϭ<���� C�a�/��� Ĉ��ЯׯC'VF�����üKG��b0��KH�K�� 
Ep�s�9���� =(�!�_�h��y�����a5�N��x��T�3lC�Ϝ�-¢�9�Kϰt�.3��}e��w�k���q'�3�JJ�͑��ϿϠ������B5P��PK�Zgt�ǿ�ߪ����߹����������$�{$�3�Z�  fUM���������Y��7�%���=�G�}�k���)Z�����  ( 5�� ������'�KY  2 E�%pIFE[@tNŰIFB�!�!� C��0� T�@į��@��*H3�� Tfx��T��T�a4��T�D=4H;
 �// */</N/`/r/�/�/�/��/�/�/�/GJ@2���5�I�v�$P�ARAM_MEN�U ?����  DEFPULS���	WAITTM�OUTT;RCV�g? SHEL�L_WRK.$CUR_STYL��;�<OPT��?�PTB�?�2C�?R?_DECSN_0<� L	OO-OVOQOcOuO �O�O�O�O�O�O�O_�._)1SSREL_�ID  ��Y��=UUSE_PRO/G %8:%*_�_>SCCRk0ORY@3��W_HOST �!8:!�T�_�ZT \Ю_ c�_�Qc<o>�[_TIMEi2OV��U)0GDEBU�GMP8;>SGINP_FLMS`�gn�hsTR�o�gPGA�`e �lC�kCH�o^�hTYPE5<A)_#_Y�}�� �������1� Z�U�g�y��������� ����	�2�-�?�Q� z�u�������ϟ��
��eWORD ?�	8;
 	PyR�`U�MAI@���SU�1E�TE�#`U��	�4R�C�OLS�n���vTR�ACECTL 1풑�B1 .I�} ~�W d�|ެ��DT Q�����РD � 7*���
��W.��.���.��`.��"���	�
��*�2�:�B�BT���"����;��3�:�B�J��+�=�O�a� s���������Ϳ߾��+Z������ ��#����������� ��;���C���K���S� ��[�����������D,�����OP��������\�nπ����Ħ �������� � �2�D�V�h�zߌ� �߰����ߦ�q�3�E� W�����ϟϱ���� _���%�7�I�[�m� ��������������� !3EWi�� 0\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z�uX�����  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲��ߚ������ 0�B�T�f�x���� ����������,�>� P�b�t����������� ����(:L^ p�������  $6HZl~ �������/  /2/D/V/h/z/�/�/ �/�/�/�/�/
??.? @?R?d?v?�?�?�?�?��?�?�?OA�$P�GTRACELE�N  A  ���@��$F_UP �����SA[@?A�T@$A_CFG ��SE=CA
T@��D�D�O�G6@��OhBDEFSPD� �sLA6@��$@H_CONF�IG �SE;C� @@dT�&3B AQP�D�Al1Q@�$@INk@?TRL �sM�A�8�EFQPE�E�W�SA�DQ�IWLIDlC�sM	�T�GRP 1�Y�b@lAC%  ���l�AA��;�H�N��R���=A!PD	� a3C	\T�Ai)iQP?� 	 �O4VGgCo ´|c^oGkB`�a�opo�o�o�o��o�b"�Bz��o7I~3 <}?�<�oN� J�����f�@)��9�_�J�`z����@
t���d�ŏ� ֏���3��W�B�{� f�x�����՟�����J�)@)
V7.10beta1�F� @�@�A&ff�QZ2�CPC�`�D��Dk`[�C�T���@ DĠ Dr[� �QBH�`�L���PC5R A?�  ��CCx����b���P!P��A����A�p�B�b!PA1������
�?L��/?333A@��"���Fff.��b�]w:�7��AeC��QKNOW_M � �E{F�TSV �Z(R�C�� ����ʿ��ٿ�$ϨA!m�SM�S�[� �B�	�E����Ϗ�̓E`
��2�E@�2���Ŵ���� L�MR�S�JY�T�j���AC5�`���e@�Rۚ]ST�Q�1 1�SK
 4	�U��A�¨߰E�� *��߽�������J� )�;�M�_�q���� ���������F�%�7�(|��Ep�2{���AG�<�����P3��������p�4��+p�5HZl~p�A6����p�7� $p�8ASe�wp�MAD0F �[Fp�OVLD  �SK�ϼOr�PARNUM  /|�O//T_SCH� [E
}'F!�)=C�%UPDF/X)�/3Tp�_CMP_O�0@T@�@'{E�$ER_CHK5yH!6
?�;RS�]��Q_M�O�o?�5_k?��__RES_GzФ~� ���?�OO�?%OO*O [ONOOrO�O�O�O�O@�O�O��3���<�? _�5��(_G_L_�3G  g_�_�_�3� �_�_�_ �3� �_o	o�3@$o CoHo�3�co�o�o�2�V 1�~կ1e��@c?��2THR_INR�0�!7³5�d�fMASS �ZwMN5sMO�N_QUEUE ��~�f��0�� *�4N0UH1NEv6;��pEND�q�?�yEcXE��u� BE�p|��sOPTIO�w��;�pPROGRAoM %hz%�p��ol/�rTASK_�I��~OCFG ��h/\���DA�TARè��@��2�����#�5�G� �k�}�������^�ן�������INFO
Ré܍�wtȟe�w� ��������ѯ���� �+�=�O�a�s����������Ϳ(�4��܌ ��I��� K_��q���T��ENB� @ͻ1>ƽ�I��G���2�� P(qO�ҡϳ� ������_EDIT �����ߋ�WE�RFL�x�cm�RG�ADJ �8�A	С�i�?�0t�
qL��q���5��?�!��<@��*�%���@�#ߊ�f�2���F�	Hp�l�G�b��>�㻎A�d�t$I��*X�/Z� **:c�0V�h���Ǟ���B��������� ����������b�� �L�B�T���x����� ����:����$, �Pb���� ���~(:h ^p������ V/ //@/6/H/�/l/ ~/�/�/�/.?�/�/? ? ?�?D?V?�?z?�? O�?�?�?�?�?rOO .O\OROdO�O�O�O�O �O�OJ_�O_4_*_<_ �_`_r_�_�_�_"o�_ �_ooo�f	���o �p�o�o�dJ��oL��o�#�oGY��PREOF ����p�p�
L�IORITY�����P�MPDS1P�>ߴwUTz�4�K�ODUCTw�e8�\�OG찇_TG;�|����rTOENT 1���� (!AF_�INE�pp�{�!�tcp{���!�ud��ˎ!�icm�����rXYڏӴ����q)�a p�/�A��p�)� j�M�Y���}������� �ן���8�J�1�n�HU�����*�s�Ӷ}}������,�?:��
jfp�/z�֯K�,�������A��,  �p�������ʿ�u"�ut�}�sF��P�PORT_NUUM�s�p�P��_CARTREP��p��|�SKSTAv�w K�LGSm���������pU�nothing�Ͽ������c{t�TEMP ����ke���_a_seiban0C�,S�y� dߝ߈��߬�����	� ���?�*�c�N��r� �����������)� �M�8�q�\�n����� ����������#I 4mX�|�������3��VE�RSI�p �d �disabl�ed>SAVE ���	260_0H721:&��!;���̏� !	(�rmoN+E/`Áeb/�/�/�/�/�*�z,�? %`���_�-� 1����E0�b8eO?a?4gnpURGE_ENB3���v�u�WF�0DO�v��vWi��4�q*��WRUP_DEL�AY �CΡ5R_HOT %�f��q:�.O�5R_NORMALH
�OrOAGSEMIQOwO�O�lqQSKIP-3���>3x$�O _1_ C_]&ot_b_�_�_�_ �_�_�_�_o(o:o o ^oLo�o�o�olo�o�o �o $�oH6X ~��h���� ���D�2�h�z������$RBTIF��4G�RCVTMO�U\�����D�CR-3��I ��QE=o�C�9.E���C���A@_�8���J]ŦU��ŉ�mĚ�n�´?[����t_V�R_ �;�x5;���0;�i;�d�u;�t�<!�A�h��R���̝�� ���&�8�J�\�n�����������RDI�O_TYPE  �4=��¯EFPO�S1 1�C�
 x/:�H2��b�M��� /��E�οi�˿ϟ� (�ÿL��pς��/� i��ϵ��ω�߭�6� ��3�l�ߐ�+ߴ�O� ���߅ߗ���2��V� ��z���9����o� ������@�R������9��������OS2 1��;+�u����-��Q���3 1�����G���>gS4 1�~����ZE~�S5 1�%7q���/�S6 1� ���/�/o/�/&/S7 1�=/O/a/��/??=?�/S8 1��/�/�/0?�?�?��?P?SMASK 1�߯ )�OF�7'XNOܯFUO_C�MOTE���X4�uA_CFG ��|M�1\A�PL_R�ANGxA���AOW_ER ���@��FSM_DRYP_RG %�%y?�!_�ETART ���N/ZUME_P�RO�O_�_X4_E�XEC_ENB � ����GSPD�dP�P�X���VTDB��_�ZRM�_�XIA_OPTIONφ�����pAINGV�ERS.a��z_�)I_AIR7PUR�@ @O�o.�=MT_�0T�@zO���OBOT_I/SOLC=N�F�1z�a�eNAMERl��bo�:OB_OR�D_NUM ?��H�aH7�21  V1wLqr�qrV0qr��sps�u\@���PC_TIME�̇��x��S232�B1����aL�TEACH PE�NDAN΀�7\H���x?c�Mai�ntenance_ ConsV2��#�"�_�No Use��N��r����������С�rNPO�>P�r\A<e�qC7H_LgP�|Nw��	<��!UD�1:b�	�R�0VA3ILRq2e��upA_SR  �:a��B�R_INT7VAL1f��I��+n��V_DATA_GRP 2��,�qs0DҐP�?`� �?��o��������կ ï�����-�/�A� w�e����������ѿ ���=�+�a�Oυ� sϕϗϩ�������� '��K�9�[߁�oߥ� ���߷���������� G�5�k�Y��}��� ���������1��U� C�e�g�y��������� ����	+Q?u�DA�$SAF_D?O_PULS�pE@p�C�� CAN�r�1f�vpSC�@��'�'Ƙ��QV0�D�D�qL�L�+AV2 y�'9K]o �������Vڈ��2($Md($C!u�1#
) @�Co/�/�/�.�W)k/ M��$�/_ @݃T:`�/�??&?39T D��3?\?n?�?�?�? �?�?�?�?�?O"O4O�FOXOjO|O֏��i%�O�O�O܉�!�L� �;�o݄��p�M
�t���Dipp�L��J� � ��jL�� �j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� ��������(�:����/c�u��� ������Ϗ��B�% �1�C�U�g�y����� ����Ƒ��0RMS �EW]�$�6�H�Z�l� ~�������Ưد��� � �2�D�V�h�z��� ����¿Կ���
�� .�@�R�d�vψϚϬ� ������M���*�<� N�`�r߄ߖߨ���� ������&�8�J�\� ǟ������������ ������,�>�P�b� p��������������� %7I[m ��������!3EWit� �OB3t����� ////A/S/e/w/�/ �/�/�/�/�*��/\?6��\R?��M	12345�678XRh!B�!̺����?�?�?�?�? �?�?OOA�>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_o] -O�_�_�_�_�_�_�_ o"o4oFoXojo|o�o8�o�oq_BH�o�o �o!3EWi{ ��������v[;�j�A�S� e�w���������я� ����+�=�O�a�xYD�k�������ɟ۟ ����#�5�G�Y�k� }�������v_ׯ��� ��1�C�U�g�y��� ������ӿ���	�ȯ -�?�Q�c�uχϙϫ� ����������)�;� M�_�σߕߧ߹��� ������%�7�I�[�@m�����v6����z��!�3�O:Cz  A�z_   �@�2�]v0� @�
��?�  	�r���`����������ph�	u�����K]o �������� #5GYk}� �0����// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-?G�p������*@  <X4�t��$SCR_G�RP 1�'�� '�� t� �t� �E5	 �1��2�2�4��W1 G3�;97�7�?�?OC���|�BD�` D��3NGK)�R-2000�iC/165F �567890���E��RC65 ��@�
1234$�E�6t�A�����C�1F�1�3�1)D�1A�:�1�I	���?_Q_c_u_�_����H��0 T�7 �2�_�?�_�_o�6�t��_Lo�_poB8bo�K�h�@�UP{��  $��1BǙ��B�  B�33Bƿ`�e�b�c�19Ag��o  @t��e�1@>@	  ?��w�bH�`2�j�1F?@ F�`\rd [o�s����� ��*��9�a�a)rU�0@�R�d�v�B���� ʏ���ُ����H� 3�l�W���{���Ě 2C�?���7����9�t�!q@"p>SԀ�D_�U�r�`y��`����G�L�3��ϯ��A>G�1��"oe$��)�t� �<�N�\�*�q�}���^� P��(����ӿ��g1EL_DEFAULT  �D���t�~��HOTSTR�� ��MIPOWE?RFL  K�ż��?�WFDO�� S�RVENT �1����P0�� L!DUM_�EIP翬��j!AF_INE�<�ϵ!FT��������!�_B� ���i�!RPC�_MAINj�Lغ8Xߵ�|�VIS��K�y����!TP�ГPU�߳�d��M�!�
PMON_PR'OXYN��e<����g��f����!RDM_SRV��r��g��1�!R�DdM���h �}�!
~��M���il���!RLSYN�@�����8��!RO�S��<�4a!�
CE�MTCO�Mb��kP�!	�vCONS���l��!vWAS�RC ���m�E!�vUSBF��n 4�0ߵ���� /�'/�K//o/��RVICE_KL� ?%�� (%�SVCPRG1�v/�*�%2�/�/� 3��/�/� 4??� 5�6?;?� 6^?c?� 7@�?�?� \��?L19�?�;�$H�O�!�/+O �!�/SO�! ?{O�!(? �O�!P?�O�!x?�O�! �?_�!�?C_�!�?k_ �!O�_�!AO�_�!iO �_�!�Oo�!�O3o�! �O[o�!	_�o�!1_�o �!Y_�o�!�_�o�!�_ {/�"� �/� F�E1 �������� 
�C�U�@�y�d����� �����Џ����?� *�c�N���r������� �̟��)��M�8� _���n�����˯��� گ�%��I�4�m�X� ��|�����ǿ�ֿ���*_DEV ~���MC:��H'�GRP 2�ׇ�+p� bx 	� 
 ,y�ϒ�+r~ϻϢ��� �������9� �]�o� Vߓ�z߷��߰����� �#�z�G���k�}�d� ������������� ��U�<�y�`����� ����*���	��- QcJ�n��� ���;"_ FX������� �/�/I/0/m/T/ �/�/�/�/�/�/�/�/ !??E?W?�{?2?�? �?�?�?�?�?O�?/O OSO:OLO�OpO�O�O �O�O�O_^?�O=_�O a_H_�_�_~_�_�_�_ �_�_o�_9oKo2ooo Vo�ozo�o�o _�o�o �o#
G.@}d �������� 1��U�<�y����o�� f�ӏ�̏	���-�?� &�c�J���n������� �ȟ����;���0� q�(���|���˯��� ֯�%��I�0�m�� f�����ǿ������R�d ��	�4���X�C�|�gϠϯ�%�x����R������ ���������+��O� =�s߁��Ϧ���i��� �������	��Q�� x��A�������� ���Y��P���)��� q�����������1� U���I��Ym� ��	�-�! E3U{i��� ���//A/// Q/w/��/�g/�/�/ �/�/??=?/d?v? -?O?)?�?�?�?�?�? OW?<O{?OoO]OO �O�O�O�O�O/O_SO �OG_5_k_Y_{_}_�_ �__�_+_�_ooCo 1ogoUowo�_�_�oo �o�o�o	?-c �o��oS�O�� ���;�}b��+� ��������ɏ�ݏ� U�:�y��m�[���� ����ş�-��Q�۟ E�3�i�W���{���� دꯡ�ï���A�/� e�S���˯���y�� ѿ����=�+�aϣ� ��ǿQϻϩ������� ���9�{�`ߟ�)ߓ� �߷ߥ�������A�g� 8�w��k�Y��}�� �������=���1��� A�g�U���y������� ���	��-=c Q������w�� �)9_�� �O����/� %/gL/^//7/// �/�/�/�/�/?/$?c/ �/W?E?g?i?{?�?�? �??�?;?�?/OOSO AOcOeOwO�O�?�OO �O_�O+__O_=___ �O�O�_�O�_�_�_o �_'ooKo�_ro�_;o �o7o�o�o�o�o�o# eoJ�o}k�� ����="�a� U�C�y�g�������ӏ ���9�Ï-��Q�?� u�c���ۏ��ҟ���� ���)��M�;�q��� ��ןa�˯��ۯݯ� %��I���p���9��� ��ǿ��׿ٿ�!�c� Hχ��{�iϟύ��� ����)�O� �_���S� A�w�eߛ߉߿���� %߯���)�O�=�s� a���߾��߇����� ��%�K�9�o���� ��_����������� !G��n��7�� ����O4F ��g���� �'/K�?/-/O/ Q/c/�/�/�/��/#/ �/??;?)?K?M?_? �?�/�?�/�?�?�?O O7O%OGO�?�?�O�? mO�O�O�O�O_�O3_ uOZ_�O#_�__�_�_ �_�_�_oM_2oq_�_ eoSo�owo�o�o�o�o %o
Io�o=+aO �s���o�!� ��9�'�]�K���� ����q���m�ۏ��� 5�#�Y�������I��� ��ßşן���1�s� X���!���y������� ��ӯ	�K�0�o���c� Q���u��������7� �G��;�)�_�Mσ� qϧ����ϗ�ߓ� �7�%�[�I���Ϧ� ��o����������3� !�W��~��G��� ��������	�/�q�V� �����w��������� ��7�.����O �s����3 �'79K�o ������#/ /3/5/G/}/��/� m/�/�/�/�/??/? �/�/|?�/U?�?�?�? �?�?�?O]?BO�?O uOO�O�O�O�O�O�O 5O_YO�OM_;_q___ �_�_�_�__�_1_�_ %ooIo7omo[o}o�o �_�o	o�o�o�o! E3i�o��Y{ U�����A�� h��1����������� ����[�@��	�s� a������������3� �W��K�9�o�]��� ��������/�ɯ#� �G�5�k�Y���ѯ�� ����{�����C� 1�gϩ���ͿW��ϯ� �������	�?߁�f� ��/ߙ߇߽߫����� ���Y�>�}��q�_� ���������� ������7�m�[���� ����������� !3iW������ }���/ e���U��� �/�/m�d/� =/�/�/�/�/�/�/? E/*?i/�/]?�/m?�? �?�?�?�??OA?�? 5O#OYOGOiO�O}O�O �?�OO�O_�O1__ U_C_e_�_�O�_�O{_ �_�_	o�_-ooQo�_ xo�oAoco=o�o�o�o �o)koP�o� q������C (�g�[�I��m��� ����ُ� �?�ɏ3� !�W�E�{�i����� ؟������/��S� A�w�����ݟg�ѯc� ����+��O���v� ��?�����Ϳ��ݿ� �'�i�Nύ�ρ�o� �ϓ��Ϸ�����A�&� e���Y�G�}�kߡߏ� ������ߵ��߱�� U�C�y�g����������$SERV_MAIL  ������OUTP�UT���RoV 2؍�  �� (����_���S�AVE���TOP�10 2�9� d 	�������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/����YP|���FZN_CFG ڍ�'��j��!?GRP 2��'&�� ,B   A�=0��D;� B�>0�  B4���RB21l�HELL�"܍�$�L��M�7�?�;%RSR�?�?�?O�?%O OIO4OmOXOjO�O�O��O�O�O�O_!_3^�  �R3_a_Xs_AR_ ��{_L�R�P�xWIR2���d�\�]�Rh6HK ;1�v; �_o "ooFooojo|o�o�o �o�o�o�o�oG�BTfb<OMM ��v?�g2FTOV_ENB��A�$���ROW_REG_�UI���IMIO/FWDL�pߥ~@5^�WAIT�r�Y��8���v@�0�T�IM�u��j�V�A��A��_UNI�T�s��$�LC�pT�RY�w$���M�ON_ALIAS� ?e�yH�he ��%�7�I�[�i���� ����m����
�� .�ٟR�d�v�����E� ��Я������*�<� N�`��q�������̿ w����&�8��\� nπϒϤ�O������� ��߻�4�F�X�j�� �ߠ߲����߁���� �0�B���f�x��� ��Y����������� >�P�b�t�������� ������(:L ��p����c� � �6HZl ~)������ / /2/D/V//z/�/ �/�/[/�/�/�/
?? �/@?R?d?v?�?3?�? �?�?�?�?�?O*O<O NO`OO�O�O�O�OeO �O�O__&_�OJ_\_ n_�_�_=_�_�_�_�_ �_�_"o4oFoXooio �o�o�o�ooo�o�o 0�oTfx�� G������,� >�P�b���������� Ώy����(�:����$SMON_D�EFPRO ����c�� *SYS�TEM*M�REC�ALL ?}c�� ( �}tp�disc 0=>�192.168.�56.1:736�0 0 ��188  Аϒ۟�����}tpconn 0 ����Пa�s�����0copy �md:picku�p.tp vir�t:\temp\���0S������/��lace��.�ӯ�d�v����7��fr�s:orderf�il.dat3�mpback>�P�ۿ�����.��b:*.*��.�ҿc�uχ�6�2x��:\,ϭ�>�0 V�������3��a�Ͻ�8���h� zߌߟ���:�U����� 
�ϸ�A���d�v�� ��,�@��������߀+߼�O�`�r����
�xyzrate 61 .�@�R�����������3700 ����dv��� ��=�<T��	�.�� �dv��� ��6�I����$� ���d/v/�/��,/ ��<V/�/�/?��/ �/> �/h?z?�?��1?@C?U?�?�?
O�#~3�13924 �? �?eOwO�O���7H @ORO�O�O_��O�O �Oa_s_�_W8�� �O?@�_�_�_$/�_ 7H�_dovo�o=,?�?@:EWo�o�oP4#? �o1N�oi{��_�_ ;oVo���o�Bo �e�w����o/A�o ��������Pa�s����? 1�?>�P�����w1�44K ՟f�x����,?�X� U����
�O��נį ֯g�y�����.�@�R� �����,���пa� sυϘ�3������ ��(���L�]�o߁�����$SNPX_�ASG 2��������7  YR%������  ?���PAR�AM ��^�� �	��P��e����*�����OFT_KB_CFG  �ô՞��OPIN_SIMW  ��%�������RVQS�TP_DSBk��%����SR ⾮� � &��OONROD��0����TOP_ON_ERR  /�W�L�PTN ����AH�RI�NG_PRMV� ���VCNT_G�P 2��'��x 	�������� ���$��VD��RP 1���(��� _q������ �%7I[m �������� /!/3/Z/W/i/{/�/ �/�/�/�/�/�/ ?? /?A?S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_r_ o_�_�_�_�_�_�_�_ �_o8o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c����������� Ϗ����)�P�M� _�q���������˟ݟ ���%�7�I�[�m� �������ܯٯ�����!�3�=PRG_�COUNTL��8�[�_�ENB��Z��M��N䑿_UPD� 1��T  
H���ۿ���(�#� 5�G�p�k�}Ϗϸϳ� ���� �����H�C� U�gߐߋߝ߯����� ���� ��-�?�h�c� u����������� ��@�;�M�_����� ������������ %7`[m�� �����83 EW�{���� ��/////X/S/ e/w/�/�/�/�/�/�/ �/?0?+?=?O?x?s?��?Q�_INFO �1�ɹ�� �F��?�?�?O�9�D��A��>>��O�3C+����BЁ@	�*7�Ң¸LY��T@P�YSDEBU)Gi�ʰ�0d��z@SP_PASSi��B?�KLOG [�ɵ���09>H�?  ����1UD1:\�D<�>�B_MPC�MɵH:_L_ɱ�Aj_ ɱ~VSAV ��M�A�A�B�5 XS�VnKTEM_TI_ME 1��G��W 0��{��rlX�O  ��T1S�VGUNSİj�'����`ASK_?OPTIONi�ɵt����?a_DI�@���[eBC2_GRP 2�ɹ�T�o�1?@�  C��cP�~�`CFG �kƧ\ b�k
}`
OB-Rxc �������� �>�)�b�M���q��� ������ˏ��(�� L�7�p����4m��� n�ϟ�\�����;� &�_�q^�QdT����� ��ѯ�������)� +�=�s�a��������� ߿Ϳ���9�'�]� Kρ�oϑϓϥ����� ������1�C���g� U�wߝߋ������߳� 	���-��Q�?�a�c� u����������� �'�M�;�q�_����� ����������7 ��Oa��!� ����!3E iW�{���� �/�///S/A/w/ e/�/�/�/�/�/�/�/ ??)?+?=?s?a?�? M�?�?�?�?O�?'O O7O]OKO�O�O�OsO �O�O�O�O_�O!_#_ 5_k_Y_�_}_�_�_�_ �_�_o�_1ooUoCo yogo�o�o�o�o�o�o �?!?Qc�o� u������� )��M�;�q�_����� ��ˏ���ݏ��7� %�G�m�[�������� ٟǟ����3�!�W� o�������ïA�� կ����A�S�e�3� ��w�����ѿ���� ��+��O�=�s�aϗ� �ϧ��ϻ������� 9�'�I�K�]ߓ߁߷� m��������#��G� 5�W�}�k������ �������1��A�C� U���y����������� ��-Q?uc ������� ��/A_q�������/� ��$TBCSG_G�RP 2���  � � 
 ?�  J/\/F/�/j/�/�/��/�/�/�/;#"*#�~1,d0?1�?!	 HD� 6s33[2�\5O1B�!x?�9�D)�6L�͞�1>���g6�0CqF�?�?�8fff�1�>��!OICj��6�1H4B�GC{OO)H��02|A�]0@HDO_O�)H�1�8CFr�O�M@  �. XU&_�O_Q_�n_9_K_�_�_�[?���0�Sp �	V�3.00�R	rwc65�S	*`��T"o�V|A�0 8 `�Y G`mHoW  � �%@�_X�o�c#!J2*#�1-��o�hCFG ���;!C!�j��B"]b�ox�BPz�Pv a������� ��<�'�`�K���o� ������ޏɏ��&� �J�5�n�Y�k����� ȟ������\	�� -�ן`�K�p������� ��ޯɯ��&�8�� \�G���k�����!/ ۿ�����5�#�Y� G�}�kϡϏϱ����� ������C�1�S�U� gߝߋ��߯�����	� ���?�-�c�Q��� Y����m������)� �M�;�q�_������� ����������%I [m9���� ���!E3i W�{����� /�///?/A/S/�/ w/�/�/�/�/�/�/? +?��C?U?g??�?�? �?�?�?�?�?OO9O KO]OoO-O�O�O�O�O �O�O�O_�O!_G_5_ k_Y_�_}_�_�_�_�_ �_o�_1ooUoCoyo go�o�o�o�o�o�o�o 	+-?uc� ���y?���� ;�)�_�M���q����� ��ݏ�����7�%� [�I��������o�ٟ ǟ����3�!�W�E� {�i���������ï�� ���A�/�e�S�u� ���������ѿ��� ��+�a��yϋϝ� G��ϻ������'�� K�9�o߁ߓߥ�c��� ��������#�5�G�� �}�k�������� ������C�1�g�U� ��y�����������	 ��-Q?a�u ������� /���q_��� ����/%/7/� /m/[/�//�/�/�/ �/�/?�/?!?3?i? W?�?{?�?�?�?�?�? O�?/OOSOAOwOeO �O�O�O�O�O�O�O_ _=_+_M_s_a_�_ C�_�_}_�_�_o9o 'o]oKo�ooo�o�o�o �o�o�o�o#Y k}�I���� �����U�C�y� g���������я��� �	�?�-�c�Q�s�u� �������ϟ��)� ;��_S�e�w�!����� ˯��ۯݯ�%��I� [�m��=�����ǿ����վ  ��� �)���$T�BJOP_GRP� 2�ݵ�  ?��i	A�H��O���� ��ߐpXd� ����� � �{,� @��`�	 �D ���CaD�q��`���fff���>��H�ϻ�L̽�	�<!a���>����=�B� � Bp��8�C�D�)�U�CQp�Dw�S�Ι��yҜ��v� ?�����?�\<���U�ҷ��%�CV+��x/���S�D5mi��{Բ��ع�<����z�>\>��33C�  CqA��`�K�j��u��bߐ���z�;�9�bB�E�>���׵ҳ� C��V���s����&��ǌ?��;��6��%�~]�D&� C����������
Ѷ� ?�s33����<Z;]u���ff�ҴK������U�)C- _i�u���� ��*IcM������Ƙ�����	V3.00�f�rc65e��* e��/ ' �F�  F��� F� F� � G� GX� G'� G;�� GR� Gj`� G�� G�|� G� G��� G�8 G��� G�< H� H� H���2 Ez  E�@� E�� EB F� FR FZ F��� F� F�P�<"G � Gp�L#?h GV� �GnH G�� �G�� G�( �=u=+*�(�$`Q�?�2�3?� � ��M?[:A��*�SYSTEM
!V�8.30218 ��38/1/201�7 A y  �p7M�TP_T�HR_TABLE�   $ $�1ENB��$D�I_NO��$D�O�4  ��1C�FG_T  �0�0MAX_IO�_SCAN�2MI�N�2_TI�2DM�E\��0@�0 � � $CO�MMENT �$CVAL	CT~�0PT_IDX��uEBL�0NUMQB�ENDIJfAZITI�D]B $DU�MMY13��$�PS_OVERF�LOW�$�F��0FLA�0YPE��2�BNC$GLB_TM�7�EF@�1�0ORQCTRL�1��$DEBU�G�CRP�@2@ � $SBR_P�AM21_VP� T$SV_ER�R_MODU4SC�L�@RACTIO��2�0GL_VIE�W�0 4 ]$PA$YtRZtR�WSPtR�A$C�A@A�6aQUeU� �0N�P3@$�GIF3@}$eQ �lP_S�PiQ L�pP�VI<P�PF�RE��VNEARPLA�N�A$F	iDI�STANCb��JOG_RADiQ�@$JOIN�TSP尤TMS�ETiQ  �WE<�UACONS2@B��RONFiQ	�? $MOU1A`��$LOCK_F�OL�A�2BGLV�@CGL�hTEST�_XM@@raEMP�E`,R�b�B`�$cUS;AfPH`2Pt�S�a�bMP_�`z�aQCENEdR~r $KARE�@}M�3TPDRAhP|;t2aVECLE�3�2dIU�aqHE�`TOOLH`�0qs�VI{sRESpIS�32�y64�3ACiHX`�`~qONLE��D29�B�pI�1�  @$RAI�L_BOXEHa�PROBO�d?�~QHOWWAR�0x�r�@�qROLM�B2�A�C �SK�r�@n�0O_F9�!��S�qiQ
>o �R�VpOCiQ_�SLiOGaK��VOUZb�R�eAELE�CTE<P`�$P{IP�fNODE�r,�r�qIN�q2^��p?CORDED�`�`�}��0P9P@ � D �@OBAU`TA�a����C�@����P�q0��ADR�A�0F@TCHup o ,�0EN�2*�1A�a_�Tl�Z@��B�RVWVA!A � ApeR�5PREV_RT�1�$EDIT��VSHWR9�S@	UА�IS`yQ$IN�D0@1QB蓗q$HEAD�5@ ��p�5@��KEyQ�@CPwSPD�JMP�yL�5�0RACE�4��a�It0S~�CHANNEzp<�	WTICK{s�1�M`A�0@�HN�AED0^�]D�`CG�qP���v�0STYf��qLO�A�3B���jP_ t 
��Gr�S%$���T=PS�?!$UNIGa5Ax�E�0�FPORT���SQU5ptR���B��TERCJ@*b�{TSG� �P�P6�$�DE��$`T�hq�0OK@>CV�IZh�D�Q�E�APR�0�AͲ�1��PU}aݵg_DObk�XSV`�K�6AXI��7��qUR_s�E$T��p��*��0FREQY_hp<�ET=�P�b��PARA`@.P
t@�[���ATHr��3@�D�s�s�0 ��2SR_Q�0ql}��@�1TRQIc0��$`�@��BRup���VE@@��NOLD���Ap7a��x@�A>��AV_MG���P��/���/�D)�D;�}DM�J_ACC.��C��<�CM��0CYaCM@3@��M@_E������٘@NbSS}C�@  hPcDS���1�@SP�0*�AT:����@��i�~�BADDRES{s=B��SHIF}b�a�_2CH�@&�I\�@|��TV�bI�2A]��h>��C�
�j�
.a����0 \��������웱�@��CnӞ�aºꯆ:R����TXSCREE���0�TIN!AWS�P;��T00r�sQ_>�jP TQ� 7P�B�6QP��
���
���RROR_�"a�@���D�1UE�G� ���U��@S�XQ�RSM�� �U�NEXg��6��0S_�S��	0���>�C�b��o� 2m6�UE���2�GRUͰGMTN_KFLQ�#POHg/BBL_�pWg@�0� ����O�QƾLEn���pTO�`C�RIGH�B�RDITd�CKGRg@�TEX,���WIDTH�sݐBh�A�A{q��I_/@�H��  8 $LT_ �|�Y0@RyP�b�s�w�B��RGOu��0D0TW�� U� �R�b�L�UM�!�^�ERV���]PFP`>��1z'@r�GEUR�ciF\��Q)��LP�Z�Ed��)'�$(P�$(�p#)5!+6!+7!+8"b�>CȰ`���F�q�aS�@�EUSReT  <��/@U�R��R�FOChq�PPRI�z�m�@?A� TRI}P�qm�UN�0
�4!�P ��0�5�p7��b;�5� "T\� ̱G �T7����}�O2OSNAd6R A���;3wq�1#n_�S �^�2�����aU!"A�$�?�?+"��;3OSFF�` P%O��3=O@ 1#PD:,D$PGUN#K`}S�B_SUBB�Pk SRT�0��&0��"avp��OR�p�E'RAU���DT�Ib���VCC��H�' ���C36MFB�1ĢSPG?�(s (b`�STE�Qaʀ9PWTѠPE�:��GXd) ����J�MOVE��{Q6RA�N4`?[�3DV�S6RLIM_X�3qV�3qV \XvQk\:V1�IP&�2VF��C砽@d��G�*��IB�P,�S� _�`�p�b����@ (0G�B�� "P�@��pr+�x �r �,� tRn@��s C@TeGDRI�PSfQV!��wdԐ��D�$MY_UBY�$\d�;QA��S���h�q�bP_�S�ף�bL�BMvkQ$j�DEYg��EX� ���BUM_�MU6�X�D<q U�S�?��;VGo�PACI�TP�<Uyr��3yrkSyr:;qRE0nr�1l�9cyrz�@,�BTARGP!P�p�R<aR{0�@�- d��;cB	4:r��R�DSWqp�S�n�:s˰O�!d�A(v�3���E��U�p0Xm�j�:cHK�.���K�AQ��0���?SE9A����WOR�@3���uMRCVr/ U��O��M�@C��	ÂC�sÂREF ��̆��gRj�
��  Ȋ�ي��=�̆r�_RC��s�����@`����b����b�to0 �Т�;��4� �e�OU���rH��\c(`+�u��2��0<���̰� -=��Ѻf�K�SUL3a.2�C7Po/+p�NT�a��]��ag��g��!g�&�L�c���cP������!�@T���s�1���o@APg_HUR�ۥSA>SCMP��F����
�_&�R�T�����X.���VGFS��E2d �M8� � Y0UF_�����J��RO� ���l�W,rUR�GR�mq�I���D_V_h[�D�@zY��3�WIN".rH���X-V
A�RqR�P�WEw�w�q`|c6v,q��RvLOiP�tc�PMc��3t� +=�PA' =�CACH6�����@��,p��2K�ۓC�Q-Io�FR"�T� $�N��$HO�@�R�� `�rc��[�֘p���ڔ�VP�r����_'SZ3p���6����12� ��]p�؆P�؛WA3�MP��aIkMGx���AD鞨qIMREٔ6�_SIZ�P��!po��6vASYNBUF6vVRTDh�t�F�~OLE_2D�T(��t��0C0aUs��yQP�X�ECCU�x�VEM�p����#�V�IRC��VTP �����G�p��t��LA�s�!���Mco�4��;�CKLA�SQC	��ђ�@5 ! �A�� @&B�Tq$��$`��6 |F@o���Xñ�T�o�?a��"�uI���r/��`�BG� VEJ�`P�K|p1���֖K�MH�O+��R7 � �}F���ESLO�W}w]RO>SAC�CE*@-�=�xVR`:��11�yrAD��/0rPA��&�D:�1�M_Ba�81N��JMP���A8y�>b�$SSC6u�2C���C��@92���S8��N/�pL;EX��: T〲Cr�Q��6�FLD?1DEZ�FIQ rO�pqty��BVP2�Ɵ;� ϱPV|多�MV_PIZ��G�BP��`а�F	IQ�PZ�$��`�����GA%�p�LOO0Tp�JC�BT*����� ��ړP�LAN�R&�L�F@���cDV�'M�p���U�$�S�P.q�% �!�%#�㱶C4G�9���RKE�1�VANC]K�A0p� <�@�?�?:Q3A�a =�?q?�?T0�9����r> hܰ�	��K9�fA2b�<X@̠OUe�ݒA���
O���SK(�M��VIE�p2= �S0:�|R? <�{@X���`UMMYR����Re��D����ACU�`b�U��@@ $�@TI}T 1$PR8��UOPT�VS�HIFʀ�A�`�a���D�0����-$�_R$�UړQ .qZ�U�s�ot�Q�av�Q5fSTG@cVSsCO��vQCNT�� �3� }w�RlW�RzV�R��W�R�XLo^opjjA2���51D>a�0�� �pSMO��B�%TC�J�@1u����_���@C%�G�i�LI� ��'��XKVR�DDY�@T��� ZABCP�E��r�b���
��ZIeP�EF%��LV���L����AZMPkCF�eGy�$p�	�rDMY_L�N$@Ar8��dH ����g��>�MCM�İC��CART_�Xq�P�1 $JvsptD��|r�r��w���u���UXW|�puUXEUL�x�q�u�t�u�q�q�y��q�v r�eI PHk�d���Y�`D�� J 8o�	V��EIGH��H?(�"��f��ĔK a�= �C���`$B&��K���1_�B��LgR�V� F�`��COVC؀qrfq9��@}�e��
����7�D�T�RȰ	�V�1�SPH� ǑL !�S�i��{����ST�S  �����_   ��� v��<�ѐNa1 ���� ������������������������	���
�����������������( ��RDI������ğ֟����t�O|����� ����ίஔ�Sz��� >�����ſ׿��� ��1�C�U�g�yϋ� �ϯ����������v� }���8�!�3�E�W�� �'�9�K�]����[ ����UЅ�� ��( ��� ��@A�v�^`BF_TT��ի����I�V>0n�J�_��I�R 1&� C8����%к� ��C�  ��������� ���"�4�F�X�j�|� ������������1 gBTjx�����р���8�0B QI�Z lJ������� ��/"/4/F/X/F� ��t/�/b*���/�/��ԋbv�@`�v�MI__CHANU� `� #3�dV�`哑&0�ET>�AD ?*��y0�m��/�/��?�?�d0RLPs��!&�!�4�?�<SNMASKn8��1_255.4E0�3�3OEOWO�OOLO�FS^Q �`�$X9O�RQCTRL �&�V�m��O��T �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo(l�OKo:ooo��;PE�pTAIL8�J�PGL_CONF�IG 	����/cell/�$CID$/grp1so�o�o1�#��?\n��� �E����"�4� �X�j�|�������A� S������0�B�я f�x���������O�� ����,�>�͟ߟt�@��������ίB�}c� ��(�:�L�^���`o��e��b���Ϳ߿� ��\�9�K�]�oρ� ��"Ϸ���������� #߲�G�Y�k�}ߏߡ� 0������������ C�U�g�y����>� ������	��-���Q� c�u�������:����� ��);��_q ����H�� %7�[m����]`�U�ser View� �i}}1234?567890�
/ /./@/R/Z$� �cz/���2�W�/�/��/�/??u/�/�3 �/d?v?�?�?�?�??�?�.4S?O*O<ONO `OrO�?�O�.5O�O �O�O__&_�OG_�.6�O�_�_�_�_�_�_9_�_�.7o_4oFoXo@jo|o�o�_�o�.8#o �o�o0B�oc�ir lCamera��o�@�����NE� ,�>�P��j�|�������ď�I  �v�)� �&�8�J�\�n���� �����ڟ����"�4�[��vR9˟���� ����ȯگ�����"� m�F�X�j�|�����G� Y�I7�����"�4� F��j�|ώ�ٿ���� ������߳�Y����� Z�l�~ߐߢߴ�[��� ����G� �2�D�V�h� z�!߃unY������� ������B�T�f��� ��������������Y� "i{�0BTfx� 1����� ,>P��Y��i�� ������/,/ >/�b/t/�/�/�/�/cu9H/�/?!?3? E?W?�h?�?�?F/�?��?�?�?OO/O�j	�u0�?jO|O�O�O�O �Ok?�O�O_�?0_B_ T_f_x_�_1OCO�p�{ ._�_�_oo+o=o�O aoso�o�_�o�o�o�o �o�_�u���oOa s���Po��� <�'�9�K�]�o� PEc����͏ߏ�� ��9�K�]������� ����ɟ۟����ϻr� '�9�K�]�o���(��� ��ɯ�����#�5� G��;�ޯ������ ɿۿ���#�5π� Y�k�}Ϗϡϳ�Z��� ��J����#�5�G�Y�  �}ߏߡ����������������   ��N�`�r��������������   $�,�J�\�n����� ������������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/�t/�/�  
��(�  �B�( 	 �/�/�/�/�/? ?8?&?H?J?\?�?�?ж?�?�?�*4� �n�O1OCO��gOyO �O�O�O�O��O�O�O _VO3_E_W_i_{_�_ �O�_�_�__�_oo /oAoSo�_wo�o�o�_ �o�o�o�o`oro Oas�o���� ��8�'�9��]� o����������ۏ� ��F�#�5�G�Y�k�}� ď֏��şן���� �1�C�U���y����� ���ӯ���	��b� ?�Q�c����������� Ͽ�(�:��)�;ς� _�qσϕϧϹ� ��� ���H�%�7�I�[�m� ��ϣߵ�������� �!�3�E�ߞ�{�� �������������� d�A�S�e�������� ������*�+r� Oas������0@ �������� ��)fr�h:\tpgl\�robots\r�2000ic6_�165f.xml �`r�����0��/����/3/ E/W/i/{/�/�/�/�/ �/�/�//
?/?A?S? e?w?�?�?�?�?�?�? �??O+O=OOOaOsO �O�O�O�O�O�O�OO _'_9_K_]_o_�_�_ �_�_�_�_�__�_#o 5oGoYoko}o�o�o�o �o�o�o o�o1C Ugy����� ��o��-�?�Q�c� u���������Ϗ��:K � 88�?�� 2��.�P�R�d����� �����П���(� R�<�^���r�����ܫ��$TPGL_O�UTPUT |���� ����%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ�Пϱ�����ˠ23�45678901 ��������0�8��� ��_�q߃ߕߧ߹�Q߀������%�7���} A�i�{����I�[� ������/�A���O� w���������W����� +=����s� ����e� '9K�Y��� ��as�/#/5/ G/Y/�g/�/�/�/�/ �/o/�/??1?C?U? �/�/�?�?�?�?�?�? }?�?O-O?OQOcO�? qO�O�O�O�O�OyO֡}�_)_;_M___q_]@��_�_� ( 	 ���_�_ o�_5o#oYoGoioko }o�o�o�o�o�o�o /UCyg�� ������	�?��Ƭ�-�G�u���c� ������ߏ���`�� ,�ΏP�b�@������ ��Οp�ޟ����:� L���p���$������� ܯ�X���$�Ư�Z� l�J������ƿؿz� ����2�DϮ�0�z� ��.ϰ��Ϡ�����b� �.���R�d�B�tߚ� �����߄����� <�N��r��&��� ������Z�l�&�8��� \�n�L���������� |����� FX�� |�0����� d0� fxV �����// �>/P/�</�/�/:/��/�/�/�/?
2�$�TPOFF_LI�M [��@W����A2N_SV�#0  �T5:P_MON S�S74�@�@2�U�1STRTCHK' S�56_=2�VTCOMPAT�J8�196VWVAR� j=�8N4 K�? O�@}2�1_DEFPR�OG %�:%?CONROD�6kO��6_DISPLA�Y*0�>?BINST�_MSK  �L� {JINUSE9R�?�DLCK�L�K�QUICKMEN��O�DSCREP�S��2tps�c�D�A1P6Y52GP_�KYST�:59RACE_CFG �F�r1�4.0	D
�?��XHNL 2E�93��Q�; $B �_�_o o2oDoVoho�zj�UITEM 2��[ �%$1�23456789y0�o�e  =<�ox�o�os  !{!@�oZC�o{ �o���9K� o/��?�e���� ��#���G���+� ��O���ŏ׏Q����� ͟ߟC��g�y���� ]������������-� ��Q��u�5�G���]� ϯ!����ſ)�տ�� �q�ϕ�����3�ݿ �ϯ���%���I�[�m� ��	ߣ�c�u��ρ��� ���3���W��)�� ?���ߌ��ߧ��� ��c�S�e�w���� ��k��������+�=� O���s�EW��c ������9� o��n��� ��#�G�"/} =/�M/s/�/��// /1/�/U/?'?9?�/ ]?�/�/�/i?�??�? �?Q?�?u?�?PO�?kO �?�O�OO�O)O;O_ʐTS�R�_UJ�g  �bUJ �Q`_UI
 m_�_z_��_8ZUD1:\��\��QR_GR�P 1�k� 	 @`@o!k�oAo/oeoSo�own� �`�o�j�a�_�o�o�e?�  '9{# YG}k���� �����C�1�g�U�w���	�E��Ï~SSCB 2%[ �!�3�E��W�i�{�����\V_�CONFIG �%]�Q]_�_���O�UTPUT <%Y�����S� e�w���������ѯ� ����+�_A@�S�e� w���������ѿ��� ��+�<�O�a�sυ� �ϩϻ��������� '�8�K�]�o߁ߓߥ� �����������#�5� F�Y�k�}������ ��������1�B�U� g�y������������� ��	->�Qcu ������� );L_q�� �����//%/ 7/H[/m//�/�/�/ �/�/�/�/?!?3?D/ W?i?{?�?�?�?�?�? �?�?OO/OAOݟ� >�O�O�O�O�O�O�O �O_!_3_E_W_J?{_ �_�_�_�_�_�_�_o o/oAoSod_wo�o�o �o�o�o�o�o+ =Oaro���� �����'�9�K� ]�n��������ɏۏ ����#�5�G�Y�j� }�������şן��� ��1�C�U�g�x��� ������ӯ���	�� -�?�Q�c�t������� ��Ͽ����)�;� M�_�p��ϕϧϹ��� ������%�7�I�[� m�~ϑߣߵ������� ���!�3�E�W�i�LH������� s���hO������1� C�U�g�y��������� t�����	-?Q cu������� �);M_q �������/ /%/7/I/[/m//�/ �/�/�/��/�/?!? 3?E?W?i?{?�?�?�? �?�?�/�?OO/OAO SOeOwO�O�O�O�O�O �?�O__+_=_O_a_ s_�_�_�_�_�_�O�_ oo'o9oKo]ooo�o �o�o�o�o�o�_�o #5GYk}�� ����o���1� C�U�g�y����������ӏ���$TX_S�CREEN 1������}��&�8�J�\�n���������ҟ� ��������P�b�t� ������!�ίE��� �(�:�L�ïp�篔� ����ʿܿ�e�w�$� 6�H�Z�l�~������ ��������� ߗ�D� ��h�zߌߞ߰���9� K���
��.�@�R��� v��ߚ����������k���$UALR�M_MSG ?��� ��zJ� \��������������� ����/"SFw+��SEV  �E���)�ECFG ���  }�u@�  A��   B��t
 x�s�0B Tfx�����~�GRP 2�w 0�v	 ��/+�I_BBL_NOTE �
�T��l��r��q� +"DE�FPRO5�%9� (%k�/�p�/�/ �/�/�/?�/%??6?�[?F??j?�?!,INUSER  o-�/�?I_MENH�IST 18�� � (|  ���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1�?`OrO�O�O��)'O9N381,2A3�O�O�O	_�O+�O�9EeditEBCONRODMOi_{_�_�_&O�O138,2��_�_�_o"o�_�_,166X_no�o�o�o�@-7oA_SR2,1�^o�o
'o�o;N4@]ov����@'?Q~2LO�
��.�Q# �0"A�?_�q������� ���CN������+� =�̏a�s��������� J�ߟ���'�9�ȟ ڟo���������ɯX� ����#�5�G�֯k� }�������ſT�f��� ��1�C�U�@�yϋ� �ϯ��������	�� -�?�Q�c��χߙ߫� ������p���)�;� M�_�q� ������ ����~��%�7�I�[� m�������������� ����!3EWi{ fϟ����� /ASew� �����/�+/ =/O/a/s/�/�/&/�/ �/�/�/??�/9?K? ]?o?�?�?"?�?�?�? �?�?O#O�?GOYOkO }O�O�O�:O�O�O�O __1_4OU_g_y_�_ �_�_>_�_�_�_	oo -o�_�_couo�o�o�o �oLo�o�o); �o_q����H Z���%�7�I���m��������Ǐ�J��$UI_PANE�DATA 1�������  	�}/�frh/cgtp�/wholedev.stmӏ1�C��U�g�R�)pri���]�}��Ɵ؟���� � )"�F�-� j�Q�������į��� �����B�T�;�x��V���  �   rP����ǿٿ���� b�3Ϧ�W�i�{ύϟ� ������������/� A�(�e�L߉ߛ߂߿�@�������� �� 8���T�Y�k�}��� �����J�����1� C�U���y���r����� ������	��-Q cJ�n��0�B� �);M�q �������/ h%//I/0/m//f/ �/�/�/�/�/�/�/!? 3??W?���?�?�? �?�?�?:?OO�AO SOeOwO�O�OO�O�O �O�O�O_ _=_O_6_ s_Z_�_�_�_�_�_�_ d?v?4O9oKo]ooo�o �o�_�o*O�o�o�o #5�oYkR�v �������1� C�*�g�N�����o"o ӏ���	��-���Q� �ou���������ϟ� H���)��M�_�F� ��j�������ݯį� ���7�����m���� ����ǿ����p�!� 3�E�W�i�{�⿟φ� ���ϼ������/�� S�:�w߉�p߭ߔ���D�V�}����-�?�Q�c�u�)	��ŉ� ��������� ���D� +�h�O�a��������� ������@R9�v	�`�Z��$UI�_POSTYPE�  `�� 	 ����QUICKMEN  ���� �RESTORE �1 `� � �i�S`N�m~�� ����/%/7/I/ [/�/�/�/�/�/r �/�/�/j/3?E?W?i? {??�?�?�?�?�?�? �?O/OAOSOeO?rO �O�OO�O�O�O__ �O=_O_a_s_�_(_�_ �_�_�_�_�O�_o"o �_Fooo�o�o�o�oZo �o�o�o#�oGY k}�:o���2 ���1�C��g�y� ��������d����	�x�-��SCRE� �?�u1�scHu2h�3�h�4h�5h�6h�7�h�8h��USER�J�O�a�TI�j�ksTr�є4є5є6є�7є8ё� NDO_CFG !�����Ѩ PDATE� ���N�one _� ��_INFO 1"`�]�0%3�x�	� f�����˯ݯ���� ��7��[�m�P��������ǿ�J�OFFS_ET %�Կ σA֏�*�<�N�{� rτϱϨϺ�Ͼ�� ��A�8�J�w�n߀�������
�����UFRAME  �ʄ�G�RTO?L_ABRT&���>�ENBG�8�GR�P 1&<Cz  A����� �������������:�� Ug��V�MS�K  j�]�X�N#���]�%�߫��oVCCM�'�V��RG��*�	���ʄƉD � BeH)�p<2C�)��PN?�` ��MR��20��p���"��р	 ���~XC56 *����Y��N�5р��A@<C� 	���ʈ); h�c��R�р|�Ђ B����6�t /T1/ /U/@/y/d/ �/�/�/�/*/�/	?�/�???�c?u?��TCC��1��f�9�рuр��GFS��22w Й�2�345678901�?�2ʈ"�6��?!O@с>,12�QO_GB@�R 8N:�o=L������ �����OOA�O�O@O _dOvO�O�O�O�_�O �O�___�_<_N_`_ r_Soeo�_Ro�o�_�_�oo&o8o��4SEGLECF�j��$�VIRTSYN�C� ��6�BqSIONTMOU-t�р��cu��3�U��U�(��� FR:\�es\+�A\�o ��� MC�vL�OG�   U�D1�vEX�с'� B@ �����q  ESK�TOP-8U37T7F�6�!�N�`��3��  =	 �1- n6  G-��ʆ�xf,p�<#�0=��ʹ����r�xTRAIAN��2�1.��
. �d��sq4w (,1��0��)�;�M� _�q���������˟ݟ����I��crSTAT 5��� ������'$��ۯ��_GE��6w�M`. �
��. 2��HOMIN��7U��U� �r(�a�a�aCG�um��JMPERR 2=8w
  �oE: ��suTs�����߿� ��'�9�O�]ώρϴ��_v_�pRE��9\t���LEX��:w�A1-e�VMPHASE  RurCCb��OFFLp�c�<vP2�t;4�0R4��8���b@�����ab>?s33��Á�1��L��ҕ�P��|��t�>x��Â���C{ASDE��R-��o��E�B��-q
.?O�W�  �E�4�B��2ҠƘ� ��� �^����<�1�`� ���`�r��� ����>����L� >��Jtn����� � �$6�&4 F\������ �j//0/Z/� �\/��/�/��/T/ �/ ??d/Y?�/z?�/ �?�/�/,?�?�?�?O N?COr?�?�?�O�?`O O�O�O�O_8O�O_ nOc_u_�O�_ _�_�_ �__o4_&oX_Mo|_ �_�_~o�o�o�o�g���TD_FILTE:t�?�� ��Wp��]o$6HZl ~������ ��)�;�M�_�q�������SHIFTM�ENU 1@x�<��%����я�� 0���f�=�O���s� ����䟻�͟����P�'�	LIVE�/SNAPD�v�sfliv�b��{�ION G�yU���menu�����:�����±���A���	����b�K�c�5M���)�@�е���A�pB8��B����Ӝѝ�������m`� ;ӥ�/�M%E��u���᱁kMO��B���z���WAITDINE�ND�3���O9KN�.�OUT#�ȹSa�4�TIM�����GϮ�@����`ϱ�ϱʞ�2�RELEASE���ĳTM�����_�ACTx��Ȫ�2�_DATA C��«�%i��ߪ���RD�IS�b��$X�VR2�D��$Z�ABC_GRP �1E8�n`,@h2\��ǽZIP1�FD�� cCo������x�MPCF_G 1G8�Bn`0<o ���=�H8�<���t� 	�w�  8R�����e�����?�k���� ��5��
\��  �a ������7�����I���z��YLIND��aJ�� �f? ,(  *s��K�p����  �//+.mN/�r/ Y/k/�/��/�/�/3/ ?�/�/J?1?n?U?�/0�?�?v�C�2K8��� ��O`o�7O@~[Ol�?�Og��A�A�ASPHER/E 2LS�?�O X?�O__>_�?�Ot_ �_?�_I_/_�_�_o �_]_:oLo�_�_�o�_ �o�o�o�o#o $67�ZZ� �k�