��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�   � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d�APPI�NFOEQ/ 9�L A �!�%N/ H� �&�)�EQUIP 2�� NAMr ��'2_OVR�$VERSI3 � �PCOUPLED�� $!PP_�� CES0s!_81�s!#J3> �! �� $SOFT��T_IDk2TO�TAL_EQs �$�0�0NO�2U SPI_INDE]��5Xk2SCREE�N_(4_2SIG�E0_?q;�0PK�_FI� 	$�THKYGPAN�E�4 � DUMMY1dDDd!OE�4LA!R�!R�	� � $TIT�!$I��N �D@d�Dd �Dc@�D5�FU6�F7�F8�F9�G0�G�GJA�E�GbA�EB�G1�G �F�G1�G�2�B!SBN_C�F>"
 8F CN�V_J� ; �"�!_�CMNT�$F�LAGS]�CH�EC�8 � ELL�SETUP ރ $HO30IO��0� %�SMAC{RO�RREPR�X� D+�0��R{�T� UTOBACK�U�0 ��)DEVIC�CT	I*0�� �0�#��`B�S$INTE�RVALO#ISP�_UNI�O`_D�O>f7uiFR_F�0AIN�1���1<c�C_WAkda^�jOFF_O0N�DEL�hL� ?aA�a1b?9a�`C#?��P�1E��#s�ATB�d��MyO� �cE D �[M�c��^qRE�V�BILrw!X�I� QrR  �� OD�P�q/$NO^PM�Wp�t�r/"�w� Яu�q�r�0D`S� p E RD_�E�pCq$FSS�Bn&$CHKBD�_SE^eAG G��"$SLOT_���2=�� V�d�%���3 a_EDI�m   � ��"��PS�`(4%�$EP�1�1$O�P�0�2�a�p_O�K�UST1P_C�� ��d��U �PLACI4!�Q�4�( �raCOMM� ,0$D����0�`��EO�WBn�IGALLOW� (K�"(2�0VARa��@�2�ao�L�0OUy�C ,Kvay��PS�`��0M_O]���w�CF�t X� �GRP0��M=qN�FLI�ܓ�0UI�RE��$g"� SW�ITCHړAX_uN�PSs"CF_��G� �� WARNM�`#!�!�qPsLI�I�NST� �COR-0bFL{TRC�TRAT�P�TE�� $ACC�1a�N ��r$OcRI�o"��RT�P�_SFg�C�HG�0I��rT(א�1�I��T�I1���� x pi#�Q��HDRBQJ; C,�2'�3'�U4'�5'�6'�7'��8'�9{5CO`T <F П����#92^��LLECy�"MULTI�b�"N���1�!���0T_}R � 4F STY �"�R`�=l�)2`�p����`T |� @�&$c�Z`�pb��Pf�MO�0�TTOӰ:�Ew�EXT����pÁB���"2� ,��[0]�}Rദ�b�}�  D"}����Q���Q�kc!���^ȇ1��bÂM���P�� Ԡ8Ë� L�  ����P��`A��$J�OBn�/�i�G�TR;IG�  d�p�� ����³�7����������_M�b! et�pF� CNG AiBA� ����M��� �!���p� �q��0��aP[`��i�*�"6����0tB񉠎"J���_Rz�gC�J���$�?�Jk�D�%C�_�;������0h ��R>�t#� �������G���0NHA;NC̳$LGa���B^a��� �D��A�`��gzRɡ�!�0�p�DB�3RA�AZ�0K�ELT�Ė��PFCT&��F�0�P��SM��cI��1� % ��% ��R��a����� S��&���M` 00{o e#HK~օA^S�������If_T$�"6SW�OCSXC)�?!%�h�p)3��T�$@�ΙPANN&�AIMG_HEIGHCr·WIDI AVT��0��H F_ASqPװ��`EXP�1|���CUST��U��&��|E\�%�C1NV _�`�a���' \%1y�`OR@�c,"�0gsk��PO��LBSYI�G��aR%��`좔Pspm��0k�DBPXWORK���(��$SKP_d�`ma�"<qTRp ) ���P��0�� �0�DJ!d/��_CN��R�#� �'PAL�S�Q�d�s�DKA7WAw'�^A�@�NFZpfBDBU��*L�"!PRS�7�
�8�Q����+ [pr�$1�$Z����Li9,v?�3ʠ��-��?�4C��.�?�4EsNEy��� /�?̈3J0RE`��20�H��CuR+$L�,C,$i3
�? =KI3NE@�K!_D�I�RO�`����ȳq0vC��h �FPAÃ3u�R�PRN�B�MR���U!�u�CR[@E�WM �SIGN���A� .q�E�Q�-$P��.$PLp 2�/ P7�PT2�PDu`L���VD�BAR@�GO_AW����Jp � �D�CS�pZ�CY_ 1���@1<�Q?fWIG2�Z2>fN>������
�qS&c}P2 oP $��RB?��e�P=hPwg�QBY�l�`gT+1�THN�DG�23��KS�SE8|�Q��SBL㸣\cc�TT.SqSL�4 HpZ ���V�TOFB�l�FE@fA�ǿb�TqSW5�b�DOC���MCS@�f�`Z$r�b H� �W0��T�!sQSL�AV�16�rIN�P��f��LyqQP�7/� $,�S����=��v��uFI��r줭sc�!��r!W1ԭrNTV'�r�rV	��uSKIvTE�@W���:��J_� _�00�S�AFE�A�_SV>��EXCLU��B ��PDJ L1�k�Yp�d�ƻrI_V� !PPLY 0b���sDE~w��_ML2��B $VRFY_4�#��Mk�IOU�� 憻 0���:�O�P��cLS�@jb;�3572$��Sr�� Px%X��{P�hs� �� 8� @� TA� qঠy � pR_SGN��96����@�A������iPt!��s"��~UN�0jdՔ�U���B �@� ��� ����KѴW I�2: @b�`Fؒ���OT�@ @�:41(�774C2�-Mv`NI�2;�R������A�q��DAY1#LOAD�T/4~��;30� �EF�X�I�b< @%1O���3� _RTRQ���= D�`@��Q.@  �EjP"�㥎�<�B�� 	�@ŏ�AMP��]>��a�����a�8Sq�D�U�@q���"CAB2��?A��0NSs���IDI�WRK�^��� V�WV_]���>� �DI��q�@�� /.�L_SE2�T���/�Z`�0�0��#�E_��u�4v�j��SWJ�j�  𲰂�	���=c�3OH�z�PPJ�v�IR!��B� ��w��d��B"����BAS h��� X ���V�����?C��Q��RQD�W��MS���AXx}�8�u�LIFE� �7�A1C�NJ���SՈ�H���Cs�>��C`QN"�U�f�OV� _�HE��N��SUP�hbC�"� _�Ԥ���_����[Q��Z��W����0��Tb��XZ$ `1V��Y2F�CM@T��$t@�N�p��!���9A `�P.�HE��SIZy֥�u�z�BN�pUFFI���p� �Q/40�<2�6C3��MSW9B� 8�KEYIMAG�CTM@A���A�Jr|#��OCVsIET���C ���V L�t���s?� Q	�!� :D�"pST�!x�0��� 0��Ѡ��0���EMAIL���@����c`__FAUL��EH�CCOU�p}$T�@��F< $d���eS]���ITvBUF��q���T  J���BdC�tp����#��SAVb $)�e�A� }���APi�e@U�b`_ H���	OT{BH�lc�Pր(0�
{��AX�1#�� @��_G�J�
�DYN_�� Gj�D�U/0veU��M����T8��F��ِ�A!H��(@u���C_r@�@K�D����=p�R���uDSPl �uPC�IMb ��J���U����Eƀ��IP�su��D���TH0�c���TuA�HSDI�ABSC�ts��0Vzp*} �$�#��NVW�G�#�$0� FJ�/d�jƓASC��U�ME�R��uFBCMPL��tETH�!AI��FU��DU �a�@;⠂CD�O � ����R_NOAUT.g` J��Pp2X��n4ĥPSm5C��%}5CI�.��k3|� =KH *}1Lp��Q��&�I� ��4#Q�6s��6ѡ�6P0��6���67�98�9�9�:J��8�:1J1�J1J1+J18J1�EJ1RJ1_J2mJ2T�;J2J2J2+JU28J2EJ2RJ2_J�3mJ3�:3KJ3PJ/�G8J3EJ3RJ�3_J4mB�1XT�>aLC`��F�f�F�5Q9g�5��FD�R�MT��V�C��C�wa}"C�RE�M,�FAj�OVM���eA�iTROVf�iDTm �jMX�l�IN�i���j�IN�D�`!�
xp /$DG���`opS�r9�D��`RIV)0�Qbj�GEAR�I%O0�K�bu�Nj�x��.؎��p�qj�Z_�MCM>�C�d`��U�R)2N ,{1��?g ��
 ?�p.I�?�qE���q!caU 0lbO����5P� �RIT5���UP2_ P Ѡ#TD= ��C�@���qP�J����C;�Q T��$9 O�)��OG��%E��3e&0IFI��e0�0̵���PT���FM�R2ieR 4vbY�vbLIq�� {g����f��Ŗb%_mAN~F�_F�I4�+�M;v`r}DGC{LF��DGDY��LD�q>t5[�5S�Sہk�S��M�? T�FS� l�T P�)���
�/$EX_)�@�)��1�� ��*�3b�5�b��G�!ieU �� p&2SWKO��D�EBUG�S��0�G�RY�zU�#BKUv� O1�@ O�PO8��Π0��Π�MS]�OO��S�M]�Eq�pQ`_?E V $�X�����TERM2�W<;�_`�ORIĀ6��X;�$Z �SM�_��$7�Y;�_0��TAy�Z;�.S��UPB�[� 9-��QbV$G����W$SEGźאE�LTO��$US]E0NFI�����p���`���X$UFR����q0豈�D5fh�OT1Ǵ TA_ ��C�NSTd�PA�TT!��Y�PTHJ�!B0En�K0�ART� ���������REL��&SHF�TF"�_���_SH"��M�!B0x� ��n�r��Z���OVR
#N&SHI����U�2= �AYLO$ 5I1�_�d���d�ERV�0*�} ��b ?�d��Q����A���RC
���ASYMh���WJ�apAE�����f�2�U��@d�5����D5��P#XGи!	�ORd�M�&��GR!���\��΢��^�����k�]� �E���TO�C�졳q��OP@��N z�3&1���aYO�a> RE��R�#b&O0��`�e���R]��������e$7PWRSpIM��[�sR_���VISy��r���UD�t�� ;^>�$H����__ADDR9fH$�AGa�z�s�i1R\� =_ H8�S�  ��S��C��C��CcSE�abaHSO0���` $���_aD`���PR�w�HTT� wUTH�a ({0�OBJE1u���-$9fLEP�-=�b � *g!AKB_qT��Sk�#DBGLV5#K�RL"�HIT�B�G0LO���TEM4$��b�������SS�p�4JQUE?RY_FLA��f QWYA���c���f� PU�"B�IO0 ��4G��H��HB� �IOLN~�d�/0i�C��$S�L�� PUT_&�$���Pwp��rSLA�� e�/2����ӡ��!��0IO F_AS:�f��$L��U ���#�04�#����,�HYOgN!'#� wUOP�g `  l!9f�b>$�`E&�!��P����'�!E&�"�&��1IP_MEMB~k0T h X #IPz�v��"_#0v� ���0��Oc6�1w��DSP�' $FO�CUSBGv�S_��UJhfi � 860S��JOG�W2�DIS�J7��O^��$J8�97���I6!�2�77_LA�BQ����0�8�1AP�HI�pQ�3�7D�+�J7JRA4`P�_�KEYp ��KILMON�j&`$XR =0c?WATCH_ �D�L��U1EL� �y`LB�k GpG�VP�-ffBCTR��fB5vbaLG|�l ���+h�"��LG_SIZ{Y��E
��F
 �FFD�HI�H�H��F �HM��F�@���C5V
� 5V
 5V�@5VM�5W�`AS)@S����@Nv1
��mx � ��R���4a�PÀU�Qk�LܲS�RDAU�UEA` I���R�PGH���� BOO~�ng� C-"2�ITGc�d��)&REC-jSgCRN)&DI(#S��RG����cl@�!#��b�!Sa�"Wkd!�T!#JG=M�gMNCH"�FN�2�fK�gPR�G�iUF�h	��hF�WD�hHL/ySTP�jV�hĀ�h`�h�RSgyH!�{&C��Es��!#���g�yU t�g�¬f|@6#�bG�i4�PO�JzZebEsM�w82�iEX'�TUI�eIP�c w��c���c���`�a�����s��Jg��KaNO�{�ANA"貇�V3AI�0zCL����?DCS_HI���������O����SI�)��S'��hIGN �@��C�aT����7DEV�wLL�єQ�6@BU𠔠oa@��T��$�GEM�'9nDcѢ��p�a@ЅC�!��O�S1��2��3��8Ք����q �T0v�-�絡.e�IDX����-fL�b�STm R�PY0����� p$E��C ���  ����dYa��r L*</��Q(6����6�EN 6�Օ~Kc_ s Y���P$ dKaD� �M�C�Rt �T0C�LDPm ��TRQ�LI`��e0x�f�FAL>1��_����DUA���LD������ORGe0�r���WX������Y���W�O�u � 	���uu���%Si�Tx��00�ް�S�[�RCLMC�i����{�m[�ՐM9I��O�v d�Q6��RQ�00�DSTB��Y� ��{a���AX��@�� �EXGCES�����M�
��w�@�¹�͡�����x(��_A@�ʊ l����V�K|��y \*�2��$M�BLIE��RE�QUIR����O���DEBU��L
�M{�zW�.!��B��i���N,03Ѩ�a{�R�RkHV�DCE�ƶTIN3 `!�TRSMw0p�S�N�����s�<�PST�  |nh�LOC9�RI� 9�EX��A��:���^��ODAQo%}��c$@�Q΂MF �A�_���p�C��P��SUP"� �F�X��IGG�"~ �0��MQ���v�5@� %����m ���m ����6#DATAd����E� 1L��v��IN�� t�+MDIF)?�!��H���1!� <�Q"ANSW�a!�ܑS�!D�)DAp��H3Q�$� ?�CU�@V_ >0���LO�P$�=ұ��	�L2����+��RR2I5� � ��QAX� d�$CALI��NUGt�2gRINp�<$RSW0���K�ABC�D_J2SE�����_J3v
p1S�P�@6 ��Pp�3P��\����J�h��P�O��IM��[�CSKP��$�P$�$J�Q[�Q,6%p%6%,'��_AZW�h!EL�����O�CMP��\��1X0R1T�Q�#�1�c@�FY�1��(�0�*Z�$�SMG�p����E�RJՐIN� ACߒ��5�bR��
1�_B�5�42d���14X҆>9DI~!��DH �30���$Vo�Y�$�a$� ��A��<�.A1��ň�H �$BEL�y lH�ACCEL�?��8���0IRCS_R��i��ATw��c�$PS �k�Lm�yP D��0G�Q<�FPATH�9WGD�3WG3&B��#�_� �2�@�AV���C;@�0�_MG|a$DDx�A@[b$FW(�����3�E�3�2�HDE��KPPABN.GR?OTSPEE�B��p_x�,!��DEFg���1m�$USE_���Pz�C ���YhP�0V� �YN���A{`uV�8uQMO�U�ANG�2�@OLGC�TINC~���B��D���W���ENCS����A�2��@INk�I&Be��Z��, VE�P'b23�_UI!<�9cLOWL3��pc x��UYfD�p��Y�� ��Uy�9C$0 fMOS`����MO����V�PERoCH  vcOV�$ �g9��c��\bYĄ�@�'�"_Ue@0��A&BuLcT����!ec�8\jWvrfTRK�%h�AY�shчq&B�u��s���&l��Rx�MOM|���h�ﰞ ���C��sYC���0DU���BS_BCKLSH_C&B��P�f �`}S�7��RB��Q.%CLAL��b?��p�X�t�CHKx�H�SN�PRTY����e������_~��d_U�Ml�ĉCу�ASC�Lބ PLMT�_AL�#��H�E�� ����E�H�-�0�Q#p_��hPC�a�h!H��ЯEǅCw��sXT�0�GCN_(1N�þ���SF�1�iV_RG�e�!��&B�n��CATΎSH~� (�D�V��f�'A��	� �@PA΄�R_	Pͅ�s_y�뀎v�`0x��s����JG5�6�̤�G`OG���rTORQUQP��c�y�@`�Ңb�q�@�_W�u �t�!�14��33��33�UI;�II�I�3F�`&������@VC�00���©�1��2�ÿ�¶�JRK�����~� DBL_SM�Q:O�Mm�_DL�1O�GRV:�3ĝ33ģ3��H_��Z@a�CcOSn˛ n�LN�� �˲��ĝ0��� ��e��ʽ̃��Z���f�cMY���z�TH�;.�THET0beN�K23�3Xҗ3��C�B]�CB�3C��AS���e��ѝ3��]��SB�3��h�GTS@! QC���'y��'<����$DU��;w�	��Q�����qQ�����$NE$T�I������)I7${0L�A�P�y��`�k�k�LP!Hn�W�1eW�S���� ������W��������Ɗ{0V��V��0��V���V��V��V��V*��V�V�H��栺��7�����H��H���H��H�H�OJ��O��OF	��O��UO��O��O��O��O�O��FW�}��	������SPBAL�ANCE�{�LE6��H_P�SP1���1��1��PFUL�C5\D\��:1=��!UTO_��ĥ�T1T2��22N ���2, ����q^<�(-B#�qTHpO~ �1>$�INSEG�2{a�REV�{`aDI�FquC91�('o21�dpOB!d�=��w�2��7P���LCHgWARR�2AB��~�u$MECH�ѰДQ�!��AX�qP�B��&r�~2�� 
p�"��1eROB�`�CR r�%��8��MSK_�4�� P �_OPR �1�(47Qst1�,`�*R(0)cB�(0|!IN�!�MTCOM�_C���0�  ��@0 �A$NO�REc�2�l ~27� 4�GR��%�FLA!$XY�Z_DA��LP;@DEBU�2 �0lR�0� ($mQCOD�S� �2�r� ��p$BUFIN�DX*P �2MO=R3� H%0�p �0��:@�p�QB�"�1���NF�TA�9Q#C�rG.B�� � $SIMUL���0�As�As�OBJE3�FAD�JUS�H�@AY_�I��xD�GOUTpΠ�4�p�P_FI�Q=8AT#�Y,`W �1P �PPQ+ 9�u�DjPFRI �PUT&0�RO�
`E+�Sp��OPWO��0��,@SYSBU<i� @$SOP�QB�y��ZU�[+ PRUYNn2�UPA;0D�V�"�Q�`_�@F��PP!�AB�!H��@IMA�GS�%0?�P!IMQAdIN$��Rc?RGOVRDEQ�R��@�QP�Pc�� L�_��feÂސRB�ߐ<pX�MC_E�D'@�  H�Ni Mx�bG��MY19F��#@EaSL30� �x $OVSL��SDIsPDEX Ǔ�f֓Hq�bV+��eN�a
��Pp�cwx�bw�o0�b_SET�0� @�Cr�%�9�RI�A3�
Vv_ ��bw{qnq|A-!�@� �4BT� àA�TUS�$TR�CA�@PB�sBTM$�w�qI�Q�d4F��s\�`0� D%0E�P�b�rr�E1"�qQpd��qEXE�p���a�"��tKs�Rp&0�p3UP�01�$Q `XNN�w���d���y� �PG|5�? $SUB�q�%�xq�q|sJMPWAeI$�Ps��LO ���1
 �E$RCV?FAIL_C@1�PÁR%P�0�#���Ȕx� �
�R_PL|s�DBTBá���PB3WD��0UM���IG�Q `�,�TNL ��b�ReQ�2��$�qP��@EǓ��|֒��DEFSP� � L%0� ��q_���CƓUNI�S��wĐe�R)��+�_�L
 P�q#@P�H_PK�5��2RETRIE|s�2�R�"@���FI�2� Ϙ $�@� �2��0DBGLV~�LOGSIZ�CH� ���U�"|�D?��g�_T:��!M�@C,
 #EM��R��y0>�8CHECKS�La��Po01��0�.�0R!LbNMKEQT��@�3�PV�n1� h�`ARp�� �1)P�2>�S�@O�R|sFORMAT�L�CO�`q����$Z��UX�P!r|A�PLIG�1� ; ˣSWIm �����,�G�AL_ G� $`@��B�a��CS2D�Q$E�1��J3DƸ�{ T�`PDCK�`|�!LbCO_J3�����T1׿� ��˰C_Q�` �; ��PAY��S2�u�_1|�2|�ȰJ�3�ИˈŬƗ�tQTWIA4��5��6S2MOMK@��������4��y0B׀AD���������PU��NR ��C���C�����4��` I$PI N�u�41�žӁ�:q� R~ȇ��ٯ��:�h� �a�֬��ց�1�'|1R\uSPEED G��0�؅��7浔؅ �%P7�m�F��U��؅SAM =G��7眪�؅MOV	B�  e0�� ��c2��v��� ���� ���c2nPsR�����İ$QH���IN 8�İ��?�[�6�؂A����X����GAMM��q�4$GETH1R@�SDe�mB
�OLIBR[�y�I�7$HI�0_5a@c2E`@#A@ 1LW^U@	�1a¬&o�ʱC=�n S`ރp �I_ ��pPmDòv�ñ'�����mD��	ȳ {�$�� 1��0IzpR� DT#|"c���~ LE^141�qw�a�?�|�MSWFuL�MȰSCRk�7�0��Ѻv���Z 0�P�@9@����2�cS_SAVEc_Dkd%]�NOe�C�q^�f� ��uϟ� }ɕQ��}���}*m+��9��ժ(��D�@���� �������b31�RA� Mam�7
5�#��^���}Mtա � ��YL��
A'�VAS 	BtRna`7GP�B
B@l3
A%`�GSB1W? ��2�2cЬ3oBB1M&@�;CL�8���G�b��1v���M!Lr�� �N�X0�d$W  @�ej@b�� @=�B D�BK�B�-�> �P�����ycİX �O�L�ñZ�E���uԣ[ ��OM� R/d/v/�/�/��A�j�M`��e�_��� | ��H ��jV��yV�� yP�ʗW�V��E���� IW��8�t��NTP=��PMp�QU�� � 8�TpQCOU,�Q�THQ�HOY2`H�YSa�ES��aU�E `"#�O��� �  �P�0�rUN��p�3��O$�J0� P�p^e������OOGRA�qk22�O�d^eITm�aB`/INFOI1���k��ak2��OI�b�{ (!SLEQ(� �a��`�foaS� ���� 4TpENA�BLBbpPTION�|s����Yw��1sGCuF��O�$J�,ñfb���R�x!��]ot:�OS_ED�ŀJ0� �N��@K��᪃ES NU��w�xAUT,!�uCOPY�����v�8 �MN���PR�UT�� �N�pOU��$Gcbn�l�_RGADJI1�2�3X_B0ݒ$ ����@��W��P������@㊀��EX�YCZLB��NS6u�N0άLGO�A�NY�Q_FREQZ�W`���+�p�\cLAm�"����Ì�uCRE�  c� IF�ѝcNmA��%i�_GmSTATUQPmMAIL�� 1��y�d����!��ELE�M�� �7 DxFEASIGq2��v���q!�er$�  I �`�"��ae�|I��ABUq�E�`D�V֑a�BAS��b� �[�Ub�r % $�y���RMS_TR C�ñj���Ca��ϑ���,r���C�YP	~ � 2� g� �DU�����Ԣ�0-��1��1���qDOUd�ceNrs��PR30z;p�rGRID�a�UsBARS(�TY�Hs��OTO�I1��P`_��!ƀ��l��O�@7t� � �`�@POR�cճ��.ֲSRV��)���DI. T���!���+��+�4)�5)�6J)�7)�8��aF���:q�M`$VAL�U|�%�ޡ��7t�� Cu'!�a��1�� (gpAN#��⛑R�p0� 1TOTcAL��[��PW��It�&�REGEN$�9��SX��sc0��Q����PTR��Z�$�_!S ��9дsV���t���rb�E��x�a�"�^b�p��V_H��DqA�C����S_Y4!��B<�S�AR�@2�� f�IG_S!Ec���˕_b`��#C_����w��?r��8%�b�H�SLG#�I1��p"=���4в�S�2̔DE�U0!Tf.p��TE�@���� !a�����Jv�,"��IL_M`K��z�н@TQ�P��a����2VF�C�T�P���^�Mu�V�1t�V1��2��2���3��3��4��4 ����С���1v�"IN	VIB@PN�; �!B2>2JU3>3J4>4J�I05���"���=p�MC_F`3 � L!!�r��M= I��M� �[PR�� KEEP_HNADD��!f�C�A�� !����"O�Q �I����"��?�"REM9!�ϲ^�uzU��e!HP�WD  S/BMSKG�a	!�B2B�
#COLLAB�!��2����4�o��`IT��A`��D� ,pF�LI@��$SYNT� ;,M�@C>��%пUP_DLYI1�MbDELAm ј��Y�PAD�A�� ��QSKIPE5� i��``On@NT�1� P_``�b�'�` �B]0�'���)3��)� �)O��*\��*i��*v���*���*9�J2�R‎��?sX��T%�|1�{2ܐ�|1��a��RDC�!F� ��pR�sR�PM�'R^��:b�2�RGE�p2��3d��FLG�Q�J�t�SsPC�c�UM_|0���2TH2NP��F@o0 1� � �x��p11���� l[P�E-Ds#ATWo�[�w�B�`�d@�A�p3�Bfc'HnP(�B��_D2gB�mOO��O�O�O�O�G3gB���O�O_ _2_D_ D_D4gB�g_y_�_P�_�_�_�G5gB��_@�_oo,o>o�G6gB��aoso�o�o�o�o +_D7gB��o�o�&8�G8gBǀ[m����US����\@ǡ`CN�h@�!uE��^�a @o��m�IO��ҍ�I���j�PO{WE!� W��: �1���0� �<5%Ȃ$DSB;����֒ �h CL@��S2;32s�� ��0�uy.��ICEU{�暐PEV@��PARsIT�њ�OPB ���FLOW�TR`2�҆]���CUN�=M�UXTA����INTERFAC�3�fU���CH�� t� � ˠ�E�A$����OM$��A�0נI����/�A�TN����Tо ��ߓ��EFA�� �"!�Ґ�� Hu!��� O�� &�*�� �����  2� �S�0~�`�	� �$3@B}%:B�Ŏ��_�DSP��JOG���V�h�_P�!s�OANq0%�0���K���_MIR���w�MT7��AP)�w�>@"���;AS������;A{PG7�BRKH����G �µ! ^���i��P��Ҏ���BS�OC��wN���1�6�SVGDE_�OP%�FSPD_�OVR�u �DLвӣOR޷�pN��b߶F_�����OV��CSF�<��
�F0Ƽ���UFRAF�TOd�LCHk"%�#OVϴ ��W[ ����8�Ң�͠;� ; @ BTIN����_$OFS��CK��WD���������r,���TR��T��_FD� �MB_)C �B��B��0��(�.Ѻ�SVe�Ґ琄�}#�G)�<�AM��B_��jթ߃_M@�~��ቂ��T�$CA����De����HBK�����I�O��թ���PPA��������Տթ�~��DVC_DB�� ?����A��,�X� b��X�3`���3�0�����ϱU󳠈�CAB�0��ˠ��c�� �Ow�UX��SUOBCPU�ˠS�0 �0�R����!�A�R��ł�!$HW_C@g@A��!��F��!�p�� � �$U r�|l�e�ATTRI���y�ˠCYC����C9A���FLT ��`������ALP׫�CHK�_SCT6��F_e�F_o���Ɓ�FS�J�j�CH�A�1��9I�s�8RSD_!聂��恩��_Tg�7�� �i�E)M,��0Mf�T&� �@�&�#�DIA�G��RAILACN���M�0�"��1`���L��{�PRB�MS   ��C4�z&�	��FUNC�"���RIN�0 "$0�7h�� S_��(@��`�0��`A��GCBL� u�A����DAp�a���LDܐð���d��j��TI�%��@�$CE_gRIAA��AF��P=�>#��D%T2b� C��a�;�OIp��DF_Lc�X�葶@�LML�FA��H�RDYO���RG��HZ 7����%MULSE� �����.k$JۺJ�����FAN_ALMsLV�1WRN5HARDr��Fk�2$SHADOW |�A���O2s�0N�r��J�_}���AU- R�+�TO_SBR ���3���:e�6�?�3_MPINF@{�8�4��3REG�N1DG�6CV��s
��FLW��m�DAL_N�:�����q��	����a�U��$�$Y_Bґ� u�_�z��� �/�EGe���ð�A#AR������2�Gܷ<�AXE��RO�B��RED��WRd��c�_�M��SY`���Ae�VSWWRI���FE�STՀ����d��Eg�)��D-�	{2��BUP��\V��]D��OTO�1)���ARY���R����6�נFIE���$�LINK�!GTH��R�T_RS��8�E��QXYZ��Z�5�VOFF���R��R�X�OB��,`8d����9cFI��Rg��􃻴,��_J$�F�貿S��q0kTu[6��1�w �a�"�b�CԀ+�DU�¤F7.�TUR0X#�eġQ�2X$P�ЩgFL��Pd���@p�UXZ8����� 1�)�KʠM��F9���ӓORQ���f&ZW30�B�OPd��,��t����A�tOV	E�qeBM���q^C�u dC�ujB�v�wL�wg��tAN=�Q�qD! fA�q��=�}��q�u�q����dC��"���ERϡj	�E��T�ńAs�@�UeX�0�W����AX��F� ���N�R��+��! +�� *�`*��`*��` *�Rp*�xp*�1�p*� � '�� 7�� G�� W� � g�� w�� ��� ��� ��đ��DEBU=�$8D3�h���RAB������sV��<� 
��i�fA ��-񷧴������a ���a���a��Rq��xq�J$�`D"�R9cLAB�Ob�u9�F�GROh��b=<��B_� ��AT�I`�0`����u8���1��ANDfp��@�����U���1ٷ �р�0�Q������PN�T$0M�SERV9E�y@� $%`dmAu�!9�PO��[0ЍP@�(�c�x@�  $]�TRQ�2
\��Bf��j�D"2�{�" � ?_ � l"T�Nc6ERRub�I��qVO`Z���TOQY��V�L�@)�1R�Ƅ G;�%�Q�2 o@^�T0�e�� ,7�ř���]�RA#� 2֓ d@����r� �Y@$�p�t ���OC�f�� � ��COUN�TUQ�FZN_C;FGe�� 4B�F��Tf4;�~�\� �
�xӭ�uC� ���M: �"fA��U��q: ��FA1 d�?&�X��@=����eB�A<�����AP��o@HEL�@��� 5��`B_BAS�3RSSRF �CSg�!��1
ש�2��3���4��5��6��7r��8
ל�ROO��йP�PNLdA�cAqBH�� ��ACK���INn�T��GB$Upq0� +\�_PU��,@0��OUJ�PHH����, u��TPF?WD_KAR��@&��REGĨ P�P�n]QUEJRO�p�`2r>0o1I0������P����6�QSEMг�O��� A�ST�Yk�SO: �4DI�w�E���r!_T}M7CMANRQ���PEND�t$K�EYSWITCH����� HE�`BoEATMW3PE�@CLE��]|� U���F>��S�DO_�HOMB O>�_�EF��PR>a9B�ABP�x�CO�!��#�O�V_M�b[0# IO�CM�d'eQ�[���HKxA� DH�QG��Ue2M�x����cFORCC�WAR�"ъ�O}M�@ � @r�T:#�0UHSP�@1&2&&3&&4�A�sЕO��L"�,�HU�NLO��c4j$E�Dt1  �SN�PX_AS��� �0+@ @��W1$S{IZ�1$VA��~�MULTIPL���#! A!� � $��� NS`��BS�ӂAC���&F'RIF�n�S��)�R� NF�ODBU$P���%B3=9Gşܪ�y@� x��SI���TE3s�r�cSG%L�1T�R$p&�П3xa�P�0STMT1q2�3P�@5VBW�p�4�SHOW�5��SmV��_G��� Rp�$PCi�oз��F�B�PHSP' A�v�Eo@VD�0vC��� ���A00 ޴RB% ZG/ ZG9 ZGTC ZG5XI6XI7XIU8XI9XIAXIBXI@ ZG3�[F8PZGFXH���XdI1qI1~I1��I1�I1�I1�I1��I1�I1�I1�I1��I1 Y1Y1Y2�WI2dI2qI2~I2�I2�I�`�X�IQp�X��I2�I2�I2�I2
 Y2Y2Y�p�hdIU3qI3~I3�I3�IU3�I3�I3�I3�IU3�I3�I3�I3 YU3Y3Y4WI4dIU4qI4~I4�I4�IU4�I4�I4�I4�IU4�I4�I4�I4 YU4Y4Y5�y5dIU5qI5~I5�I5�IU5�I5�I5�I5�IU5�I5�I5�I5 YU5Y5Y6�y6dIU6qI6~I6�I6�IU6�I6�I6�I6�IU6�I6�I6�I6 YU6Y6Y7�y7dIU7qI7~I7�I7�IU7�I7�I7�I7�IU7�I7�I7�I7 Ye7Y7T�VP� =Uc�� l�נ���
>A820�����RCM2���MbT�R��|���Q_�ЁR-��ń�����Y�SL�1�� � �%^2��-4�'4��x-Y�BVALU��Ё���)���FJ�ID�_L���HI��I��LE_������$OE�SAb��� h 7�VE_BLCK¡1>'�D_CPU7ɩ  7ɝ �����E����R � � �PW��>�E ��LA��1Saѝî���R?UN_FLG�Ŝ� ����� ���������šH���Ч��T�BC2��� � _ B��� br� 8W?�eTDC�����X��3f�S�TH�e�����R>�k�ESERVEX��e®�3�2 �d��� ��X -$��L�ENX��e�Ѕ�RyA��3�LOW_7��d�1��Ҵ2 �MO$/�s%S80t�I��"�`ޱH����]�DEm�41LACE�2�CqCr#"�_MA� pl��|��TCV����|�T�������0B k�)A�|�)AJ��%E�M7���J��B@k�X�|���2p �0:@�q�j�x JK��VK�X�����ы�J0l����JJ��JJ��AAL���������e4��5�Ӵ N1��P ����LF�_�1�� � �CF�"�{ `�GROU��(�1�AN6�C�#\ ?REQUIR��4�EBU�#��8�$Tm�2���|�ܑ %�� \�AP�PR� CA�
$�OPEN�CLO�S<�Sv��	k�
\��&� �<�Mh�p����v"/_MG�9CD@�C ��D�BRKBNOLD|B�0RTMO_7�H�r3J��P�� ������������6��1�@ �H!�%��� �� ���'��-#PATH)'B!8#B!��>#� � �@�1SCaA���8IN�ңUCL�]1� C2@UM�(Y"��#�"������*���*��� PAYwLOA�J2LڠOR_AN`�3L���9
1�)1CR_F�2LSHi2D4LO�4�!H7�#V7�#ACRL_�%�0�'�$r��H���$HC^�2FLEX�;J#�� P�4�F�Э߿�2��J��� :����|�HG_D�����|���'�F1 _A�E�G6�H�Z�l�~����BE�������� ����*��X�T,�C� ���@�XK�]�o�^Av�	T&g�QX>�?��4T X���eoX�������� ����������	-	:�J@� �/�M0_q~�۠AT�F��6�ELHP���s�Jڗ � JEoCTR�!�ATN���v|HAND_VB�q�1��$� $:`�F2Cx���SW��"�� $$M,00�_Y�n i��P\����A��� 3����<AM��_AmA|��NP�_UDmD|P\ G���E�STaM�nM�NDY��� C���� 0��>7_A>7Y1�'��d�@i`�P���@����""J$�� O�4D'"r�J�<��ASYMl%A�	� l&��@�-Y1�/_�}8� �$��� � �/�/�/�/3J	<��:;�1�:9�D_VI��x���V_UCNI�ӝ��cF1J�� ��䕶�Y<��p5Ǵ� y=6��9��?�?>�wc��4�3��$�� ASS  ���s�=� |�h�VERSIONp�w �
���IRTU<�qσ�A�AVM_WRK �2 ��� 0  �5�z�������� �	8�)�L�=�B���:�w�^�|�(� �ݧ�7ѭ����������BSPOS� 1���� <��A�S�e�w��� �����������+� =�O�a�s��������� ������'9K ]o������ ��#5GYk }��������//1/C/U/ⰑA�XLMT��X#�n%�  dj$INs/��!i$PRE_EXE�(� �&)0�q��������LARMRECOV ����"
�LMDG �����[/LM_IF �ˆ!X/ c?u?�?�?�:Q?�?�?x�? OM, 
0� 8O�4�cOuO�O�O��NGTOL  <���A   �O�K���PP)�O ; ?6_,_>_P_{� $BR_�_w�o_ �_�_�_�_�_o�_'oo7o]o�!��O�o�o �o�o�o�o�o+�=Oa�PPLI7CAT��?��� ��J`Ha�ndlingTo�ol �u 
V�8.30P/33��@lt��
8�8340�slu

F0�q�z=�?
2026�tlu���_��7DC3�pJ � �sNonelx� FRA�߇����B�T�IV�%�s�#��U_TOMOD� E��)P_CHGAP�ON������ҀOUPLED 1��� ��"�4�uz�_CUREQ 1M��  � >�>��*ސ�4��!��x�{~� ��uƄ�Hm����HTTHKY����w� ��7����%�C�I�[� m��������ǯٯ3� ���!�?�E�W�i�{� ������ÿտ/���� �;�A�S�e�wωϛ� �Ͽ���+�����7� =�O�a�s߅ߗߩ߻� ��'�����3�9�K� ]�o�������#� �����/�5�G�Y�k� }������������� +1CUgy� �����	' -?Qcu��� �/��/#/)/;/ M/_/q/�/�/�/�/? �/�/??%?7?I?[?0m??��P�TO�@�����DO_CLEA�N܏��CNM  �K >�aOsO��O�O�OD�DSPDgRYRO̅HI��=M@NO_'_9_K_]_ o_�_�_�_�_�_�_�_J�MAX�p�4�1���aX�4"��"���PLUGG���7����PRC�@B;@"?K_�_ebOjb�O^��SEGFӀK�o �g�a;OMO'9K8]�o�aLAP�O~ Ǔ��������/�A�S�e�w���΃T�OTAL-fVi΃U�SENU�`�� �䏺�P�RGDI_SPMMC�`{q�C�aa@@}r��O��@f�e��_STRING 1	ˋ�
�MĀS���
`�_ITE;M1j�  n���� ������Ο����� (�:�L�^�p����������ʯܯI/O SIGNALd��Tryout� Modek�I�np�Simul�atedo�Ou�t.�OVER�R�@ = 100�n�In cyc�l"�o�Prog� Abor8�o�~�Statusm��	Heartbe�ati�MH F�aul����Aler���ݿ���%��7�I�[�m��  �3f��1x��������� ��*�<�N�`�r߄� �ߨߺ�����������WOR�`f�L��� &�t��������� ����(�:�L�^�p������������PO d�����d���%7 I[m���� ���!3EWi��DEV��� �����//'/ 9/K/]/o/�/�/�/�/��/�/�/�/?PALT��81d�?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O�O&?GRI`f��A P?�O__(_:_L_^_ p_�_�_�_�_�_�_�_� oo$o6oHo�OR �̀a�OZo�o�o�o�o �o&8J\n �������noPREG<>%��o� L�^�p���������ʏ ܏� ��$�6�H�Z��l�~�����$AR�G_L�D ?	����ӑ��  	$��	[�]�����ƐSBN_C�ONFIG 
�ӛ&�%� �CI�I_SAVE  ��E�<�ƐTC�ELLSETUP� Ӛ%  O�ME_IO��%?MOV_H�������REP�l���U�TOBACKt��0�FRA:\�� ���_�'�`���=�� J� 	�������ͿĿֿ�6����	�1�C�U�g�yϋ� �Ϸ���������� ��5�G�Y�k�}ߏߡ� ,������������ C�U�g�y����aׁ  )�_�_\�ATBCKCTL�.TMP DATE.D;<��	��-�\?��INI;0p��8��MESSA�GT�^�_�ېi�ODE_D��W�8�H����O����PAUS���!�ӛ ((O֒��
��* N<r`��������"����TSK  ��=�C��	�UPDT��\�d����XWZD_�ENB\�4��ST�A[�ӑ�őXIS~&�UNT 2ӕ�`� � 	S���c2�V�0�D�[* Qs����  �`	'$h�
/L/^. "�YK����J'"��b}�2c/�/_/�/�/��MET�`2�P�/?�/<?�)SCR�DCFG 1C/`��\�\�1?�?�?�?�?�?�?6��QX��??OQOcO uO�O�O O�O$O�O�O __)_;_�O�O����GR����zS��N5A��қ	�wV�_EDZ�1e9��9 �%-��ED�T-h_ʪ�_o�`/�A���-��_��	������_�o  ���e2�oɫko�o �6k�o!hozo�o�c3Y�o��o�n�@�4F�j�c4%� �r���nN��� ����6��c5�a�>��� �n���̏ޏt���c6��-�
�Q��n�Q� ����@�Ο�c7���� ֯��n���d�v������c8U��_����0
 }~��0�B�ؿf�B�c9!ϑ�nϵ� }�Jϵ���Ϥ�2φaCR�oį9�K����������n���zP�PNO�_DEL�_xRGE?_UNUSE�_vT�IGALLOW �1�Y~�(�*SYSTEM*� 3	$SERV�_GR�R 69���REGB�$d� <9��NUMg��z�P�MU�� 5LA�Y�  <PM�PAL[��CYC10����������ULSU��{������D�L�N�BOX�ORIk�CUR_�;�z�PMCNV6��;�10���T4DLI�4�V����ߨ��'�9K]oR�zPLA�L_OUT �Dcc�QWD_AB�OR��	��ITR/_RTN���Y� �NONS8� ��CE_RIA_UI��<F_1���B =[_�PARAMGP �1�w�`_����Cp U .� � � U� � � � U� � � � �� �  D5`DQ$3!g-�<$�H$}�T$� DX �� X "� B�D�1� 9X @� 6?� <HE��ONFqIy���!G_P��;1� �e�U ??0?B?T?f?x?�?��!KPAUSX�19�UR ,Z��? �?�?�?�?OOOTO >OxObO�O�O�O�O�Oh�O_�2O_e�y�PCOLLECT__�Y5auGW�EN��I�"cR QN[DEOS�W����1234567890�W�S�u8�_�Vy
 H�y)�_#oS��_ohoT� AoSo�owo�o�o�o�o �o�o<+�O as������ ��\�'�9�K���o�l�VQ�2W[ � |t�VIO �YcQyH&�8�J�\���TR�2؍(Ć�
��j��  �����%�_MOR�҂!� + �'� 	 �5�#�Y�G� }�k����Ӂ"��2�?�!�!3 ҡ�KTڤ��$R_#*_�	���C4  A�S yC  x�A�3!z  BC!�PB|/!�PC  @*�����:d�U
�IPS$����T��FPROG �%�*6߼�8��I�����&RҴKEY?_TBL  )VR�� �	
��� !"#$�%&'()*+,�-./�W:;<=�>?@ABC��G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~��������������������������������������������������������������������������������͓���������������������������������耇�����������������������1��LC�Kۼ3���STA��д_AUT��Or(��U�INDtT<D�FQR_T1_�Q׃T2��7$����X�C� 2����P8�
SONY X�C-56��ྒ��@���u� ���А�HCR5��cT0�B�7T�f�Affrꬿ���� �������5�G� "�k�}�X��������������ǼTRL^��LETEG���T_SCREEN� �*kc�sc:U$MME�NU 1&�)  <���y ��Ã�= &sJ\���� ���'/�/]/4/ F/l/�/|/�/�/�/�/ ?�/�/ ?Y?0?B?�? f?x?�?�?�?�?O�? �?COO,OyOPObO�O �O�O�O�O�O�O-__ _<_u_L_^_�_�_�_ �_�_�_�_)o oo_o 6oHo�olo~o�o�o�o �o�o�oI 2X��hz���� _M�ANUAL�ߕ�D�B��L+�DBG�_ERRL��'�� �\�n�����NUMLI�MK�d �p�D�BPXWORK 1(�I�ޏ�����&�ŽDBTB_�@ )��������qDB_AW�AY�_�GCP�  �=�װ�~�_CAL��D�z��Y���M � �_)� 1*V����
͏`����6�@�_M{ГISAЉ�@B�P�OoNTIMJ� ���p�ƙ
�ۓM?OTNEND߿ڔ�RECORD 1�0}� �>�?�G�O����?���2� D�V�h���p������ *�߿�Ϛ���9Ϩ� ]�̿�ϓϥϷ�R��� J���n�#�5�G�Y��� }��ϡ���������� j���C��g�y�� �����0���T�	�� -�?���c���\���� ������P�����; ��_q�����( �L%�4[ �����^t �l!/�E/W/i/{/ /�//�/2/�/�/?�?�/z�TOLER7ENC��B�В���L���CSS_�CNSTCY 1�16�  ?Β� �?�?�?�?�?�?�?O O&O8OJO`OnO�O�O�O�O�O�Oc4DEV�ICE 126� b�*_?_Q_c_u_ �_�_�_�_�_�_?�d3�HNDGD 3�6�Cz�^LS 24]�__oqo�o��o�o�o�o�_e2PA?RAM 5�B���t�dc4SLAV�E 66�e_C�FG 7��gd�MC:\e0L�%04d.CSV��o��c|�r�"A &�sCH�p&a&��n(��w��f�r�����ÀJP��>��\_CRC_O_UT 8U�����oEpSGN 9�U�Ƣ��\��15-OCT-22 19:13�p��02��4:�41�p9V UBu1�݁�nހ���o��Im��P��uG��@uVE�RSION ���V3.5.�11E�EFLOG�IC 1:ݫ 	6��|�C����^�PROG_EN�B����͢��ULS�{� ��^�_AC�CLIM|���Xs��WRST�JN[���ţ�^�M�O��¡Zr,�INI�T ;ݪs5� �*�OPT$p ?�	i�B�
 	�R575�c��74j��6��7��50��R�Ƣ2��6��X�y�TO  ���?��Y�VP�DEX�d����@W�PATHw A��A\E������7;IAG_G�RP 2@�k�,�"	 E� � F?h Fx� E?`�D��@û��V1"�ü��T0�K�9�Cf�py�pY��dC�pq��B�i�ùm�p4m5 7890123456���;����  A��ffA�=qA�ةpхA��WHAĩp������?�A��Mk���@��tp�p��W0�A�T0T0�pB4�ü Qô���
����(�A�A��
=A�L����A��
A�Q��A�������� e�����e� Pe�:�_�{A�d������dѩp�������A����������r߄ߖߨߺ�@�EG��A@�p:�RAU5d�/��)��#P�d�l������"��4�F�@�Pz�AJ���c�?��9p�A�3\)A,��A&����0���������@�cP�]���AW�P�J��C���<d�4�-d�%G��(�:�L�^�@� ��$HZ��. |����bt�  2Vh�xm� ����[���s������=�
==�G���>�Ĝ��7���8��b��7�7�%�@�;�\"&�p�.%���@�Ah�p9 A���<i��<xn�;=R�=s���=x<�=�~�Z�;��%<�'�'�~ �?+�ƨC�  <(��U� 4"�;���&����%ùf��@?Œ?�? @?R?g��$^?�?"?�?�?�?�?�?�?)7�L?S�FB$��/"Eͽ�>OG��ΐԬq��sD�L4�x�CA��Gb�t� ����-_7_�C��_�;�/_�NED  �E�  Eh� 	D[PbRD_¿�_��8�?�����z�9�=�P�Q3�3�n������?��pDP�O=�V/�D@��<�{_�_w_o�K:o@bù��Y6�d�6`����A�U!o�o
o�o�o�o��o�oĿDICT_�CONFIG ΂�Yt؃�eg��ԱSTB_F_TTS�
ę�Vs3���
�iv[�M�AU���Y�MSW_CF*pB�s�!��OCVIEW}pC�}���6�
�� .�@�R�d�w����� ��ȏڏ�{��"�4� F�X�j���������ğ ֟������0�B�T� f�x��������ү� �����,�>�P�b�t� �������ο��� ��(�:�L�^�pς��|KRC�sDJ�r!� �κ�������7�&��[�otSBL_FA?ULT E���x>u�GPMSK_w���pTDIAG �F.y�q�IU�D1: 6789?012345��;x�MP�o!�3�E�W�i� {������������`��/�A��( W!��J�"
��vTR'ECP����
���� �M�(:L^ p�������  $6]�o�l���UMP_OPTIcON_p�ގTR�rt`s���PME^u��Y_TEMP � È�3B��pp �A  �UN�I�pau!�vYN_?BRK G�y���EMGDI_ST�A%�1!�rL NC6S#1H�{ �K��9�/_}dd�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO��O�O�O �O�I�!�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo Xo�JO�o�o�o�o�O �o�o+=Oa s������� ��'�9�K�]�wo�� �������oۏ���� #�5�G�Y�k�}����� ��şן�����1� C�U�o�]�������ɏ �����	��-�?�Q� c�u���������Ͽ� ���)�;�M�g�y� �ϕϧ�]�ӯ����� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�_�q�{���� ����������/�A� S�e�w����������� ����+=Oi� s�������� '9K]o� �������/ #/5/G/ak/}/�/�/ ��/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OY/ KOuO�O�O�/�/�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oQOcOmoo�o �o�O�o�o�o�o! 3EWi{��� ������/��o [oe�w������o��я �����+�=�O�a� s���������͟ߟ� ��'�9�S�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� K�9�g�yϋϥ����� ������	��-�?�Q� c�u߇ߙ߽߫����� ����)�C�U�_�q� ��9�Ϲ�������� �%�7�I�[�m���� ������������! ;�M�Wi{��� ����/A Sew����� ��//+/EO/a/ s/�/��/�/�/�/�/ ??'?9?K?]?o?�? �?�?�?�?�?�?�?O #O=/GOYOkO}O�/�O �O�O�O�O�O__1_ C_U_g_y_�_�_�_�_ �_�_�_	oo5O'oQo couo�O�O�o�o�o�o �o);M_q �������� �-o?oI�[�m���o ����Ǐُ����!� 3�E�W�i�{������� ß՟������7�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��/�9�K�]�oω� �ϥϷ���������� #�5�G�Y�k�}ߏߡ� �����������'�� C�U�g��w����� ������	��-�?�Q� c�u������������� ���1�;M_ ������� %7I[m� ������) 3/E/W/i/��/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�? �?�?O!/+O=OOOaO {/�O�O�O�O�O�O�O __'_9_K_]_o_�_ �_�_�_�_�_�_�_O #o5oGoYosOeo�o�o �o�o�o�o�o1 CUgy���� ���o�-�?�Q� ko}o��������Ϗ� ���)�;�M�_�q� ��������˟ݟ�	� �%�7�I�[�u���� ����ǯٯ����!� 3�E�W�i�{������� ÿտ�a���/�A� S�m�wωϛϭϿ��� ������+�=�O�a� s߅ߗߩ߻������� ��'�9�K�e�o�� ������������� #�5�G�Y�k�}����� �����������1 C]�Sy���� ���	-?Q cu��������� �$ENETMODE 1I^��    (/:+�
 RROR_PR_OG %*%�}/�)X%TABLE  +h�/�/��/�'X"SEV_N�UM &"  ��!!0X!_A�UTO_ENB � D%#U$_NON21 J+9!2_  *�u0�u0%�u0�u0(0+t0�?8�?�?N4HIS3
� G;_ALM 1]K+ �u< +�?/OAOSOeO�wO�O�?_2T0  �+s1:"�J
 T�CP_VER �!*!u/�O$EX�TLOG_REQ��6�E9 SSIZ\)_TSTKFYc5��RTOL  �
Dz�2�A= T_BWD�@�P�<6�Q8W_DI�Q L^G48$
<?"�VSTEP�_�_|
 �POP_DOh_�!FDR_GRP� 1M)B1d 	��Ofo: W`�������glp�w�qŗ���I �����fWc�o�mW`C}��XB�_�A����AX�A� ��B�;��mB��"B<A����@!�A�?zB��m�o 3WB{f���  A�PKA"?��>�Β� 
 E�� �a�q�rhN��B���8�#�\��m`}d�C��N��B�y{���m@UUT���UTF�Ϗj��s����m�OHcEP]���O��#M���*�KA���m?��F��:6:�N�r�9-��z���  �$7@��v�
�������-��+FE�ATURE N�^�P>!H�andlingT�ool � mp�BoEngl�ish Dict�ionary��
PR4D �Stڐard� � ox, A�nalog I/�O�  ct\b�+�gle Shi�ft�  !*�u�to Softw�are Upda�te  fd -�c�matic B�ackup�IF� O��gro�und Edit�ސ�g R6�Camera3�F�7�Part��nr�RndIm���p�shi��ommo�n calib �U���n����Mo�nitor�Ca�lM�tr�Re�liabL��RI�NTData Acquis��Z�ϠC�iagnoqs��0�<�almC��ocument Viewe�\����C�ual Che�ck Safet�y��  - B�E�nhanced �Us��Fr���8� R5�xt. oDIO �fin�s (�@ϲend���Err�Lm� D� p^���s	�E%N�r.�հ �P��rdsFCT�N Menu��v�8���m�FTP ;In'�facN�=��G��p Mask� Exc��gǱi�sp��HT^�Pr�oxy Sv�� � VLOAאig�h-Spe��Sk�iݤ ef.>�H�f�ٰmmunicons�
!�
��urE�'�7�r�t F4�a�c�onnect 2�;�Incr`�st�ru���� Sp�KAREL C�md. L��uaΊ�OAD*�=�Ru�n-TiưEnv�� �D;�(�el u+��s��S/W��.{�Lice'nse����
�����ogBook(S?ystem)蔭��JMACRO�s,��/OffseS�Z�MHٰp���� j73ΰMMRx��l�35.f��echStop��yt�R� ize*�3Mi��O� 2�7��x��0����miz���odM�witc�h����a�.�� yv���Optm���49���filN��ORD��0�g��� 8496�ult�i-T������C�PCM fuyn,��.sv�oO���� �^�5�/Regi��r��	��!2�ri��F� � H59k�1�Nu�m Sel*�  �74 H��İ A�dju���adi�n��O� ,[���t'atub��\У��������RDM R�obot��sco�ve� �d e�m(�ٱn� SW|��Servoٰ�s�ꒄ�SNPX b��1��g P��Libr���1�ڐ 9� ɰW.30g o��tE�ossag� f���@ e����"Lg��/I_�
�I�?TMILIB���~� P Firmn�p��^�F�Acc��x��0���TPTX����510.� el�n���������Hw573�rquM��imula��� �2�Touz�Paxѩ1� T��6����&��ev.��IUSB po�����iP�a�� 0�\sy nexc�ept��3 <� \�h51 ����oduV#��9���Q�VN�k"6PCV�L{&�^}$SP /CSUI�d���+�XC��auҠWeOb Pl���t?  �#S��\"	2��������S�&ު�V?8G�ridplay���&� ��8�-iR�b".� @ � R-�2000iC/1�65¦ d+�+�l�arm Cause/1 ed�<0:ПAscii����L�oad��V4�3Upql�0�_CycL��c�m�ori����F�RA[�am�) t{dt��NRTLi��3Onݐe He�lݨ 542*�P	C`ρ�4�`�]�1�trߵ48��RO_S Ethv�t[�ܿ�10\ҠiR�}$2D PkߵD�ER>1�E����of��A��ΰ�FIm��F��� z��64MB DRAMު�@:��9RFROA[�Ce�ll3� ����shrQ
��Zc���ÍUk�}p� pide�W�tyL�s��|0\$z�!CtdѰ�.��@"oEmai��li����+�\�� R0�q�Z$GigE�N�4OL�@Sup"��b�pW3oa�~�cro�� ����4��QM��Fauest�A>�j�� miH9.dVir�t��W��0{&Im�M�+T���}$Ko�l/ Bui��n�յ'GAPL�&��MyV6�s "�0�*CGP�Yl���{RG�'p�{�SBUW�RQ�)K�&cm\:��z��fXb�)O�võ(TA�&'spoҠ-�B�&���
 I�\E P�+�C�B'fg-��&"�  �E��sv �b��vv�3��S_k���TO;-�EH�f6.:
�E�vfx_z�)�V��tr>�)�hZ%.�F�& � ��r���*�G�&���њr�����H��РJzCTIeAc�pw4�LN�:1�Mr�" #[��Dg�"�M�-�P2��~T�@����vxuIi�-�S�&�S�&��*4�W��2.pc�)VGF��fxw�ʪVP2AU \f1x���N�if�u����"in��VPB^���)��s�D���*�a<s�F�5 �M��s�I��wc�{&Traİ���U,p  ��<���2��RDp	��N��HY���p���-��H���Øp)����� �ϭ����ħ���rдy����í4+�Ϟ�'9L���ӎ��y�9ӫ�yc3�U��B�Oߞq�u��kߍӍ�Sy*�ߩ�\Yyy����k�W�ߞ�ӄ�Yx����:��	�����y��5�o�e/�Q��,�K�m���g��^9~���u�2��A���������F�y�����y�)����|����1�m��.�+�M��8<G�i�7n��c����1�� �����W�����7�{<����6�Z�������uk��[�3|�!��?�ϔ�s�iB\����_F��{�x@.��wrst���B<�� H68���@H)T@J�EE�NDI?��tql[}
_�w�P��TQ (��IG) "���PA�p��T�/��85/A#bs;/�C/U/� ,q�/B�Gp�/�#��/�"36�5�R ?!2Oepai?5!:/pY4W���%INTo? e?_.q�?4)��?�2�pa2g�?�F �O�?A�ad6?��ty ZUD2gunOO�qC533R?�D�0u�O�/�Mcm���OO�LNT�?��P_�����0_QR7�L_�Cfi�._H?_,_f'R50<�_�SAF-F�_�7�w.vo��_�_88�/�dM Cbo����o�bvrEo��p�aa�oaD�@�osF'-AS-sS�p'�Is(�PCesXPL��O�tlo_�ut\�a�Oh%afvh%- B��/����C�$��srp�?@_�?�`w�}�bA�����h��`��]T�ˏ�sg#ch�os�t��CG\s;��us�?���sSg�/�G J��&��GDǟi$"�o�ggdiʏ!�fd��8�?h%J64S��Tut�o�O�?s����F �_����E�0���D`!�)�NO4E�O�fi$II���iwjO�l�ž��>�?*�lb
��V��vjr/��
� ��7��ϥ�_�?zG7\2O�EG��Ϲ?�`��1� ޯ��_d�o�i�8��c�50�>�x�Ͻ�"Lo�h%����dj9�﴿ƿؿ��c� up9�C� #j9{�E��L��Ek,B串����oS_�e_�&/��O}�j94JϬ�duZ��U����=d;�����8���r7�Dhu���;]m T������d��f�a����M����P�-4r 8V��O" #S�d3wc�P�in�`��a�?& HTuR�ef���
�?hcĕg�r"��q.JG	"�erM/��/ ̢/LRA^��uH7�1�/�tCK�/<eT�XP/?i�k1/m5k3.f��riR�ecHG�/�/ cr��NHGRf?L�i�Y�7�hOuX��H\m O��oρ�;H��DD@ �O��*�<�:I�?�?��8d�R�_ hd�g�hgOO�_���gm	h�_h�m��XO�o|O@�O�o�O\/�o0�f�gm�o`��`e۠;iov��yt��"���uR60���#t1mo_�#1��fdr,op7��_����lp>oh���冬~ ߏ�dLgts���&dޏ��/�o�o
�J?<�vr�F���v.R���Ɵpld�56�%4�0�/���reeK�m�X�P)�KCO*O|%56?�OZ� o~����E$io����jߠ���3l ����OR��LcOFvod��_IF��@$�� ߪ�DߦX!B�f Uce��t�4 �&��(M�O�5)e?Ƕ�/���1?Q�D�uk�'�|����`�boto�����-���6�p`�eS ��on*� ��^�lB'����Տ_�8q�_�rdk��4f ��C(ҿȿ¯ԯ�������̟�����
9I��571��t�gadi39Tar��l�ofk�������v3Pa�@� PJ��|*�������f�et�4epg��2�ed�� E�5��RI  �H552� 747��21�pWel/R78�,� ��0ETXJ6�14��ATUP  wmfh G545�p�"6�p�k�VCAM � 7\awC{RI@ ED" G �UIF)!28 { j�CNREM���`�63�a�S�CH  4C �DOCV� CS�Ui�!0 D s�EIOCE�5�4�#R694 w=e!!ESET=S#!�3!�a 73!fanuMASK��?PRXY�_"q7� �0�OCO���"3=P[�#"�ER� J�" 7�!!J�774#!39�  �Eq�G1�LCH� 0#OPLG%J�5000#MHCR�)%PS�17#MCS� 4D"�04 O#J5y5 [#MDSWe!fY1MD#1s#OP#1.#MPR$07�0w"�0�#�  �#PCMX �#R0A�#� & �00�#� ( �&0�$s50( �#PRS� �3J6903FR�D@ 02RMCNny�ndM�93 ~SNBAA��800�@HLB o "Lo�SM�A�0 (Ww"4 on�it#!2  II�)�TC [#TM�ILe �B�`0"K3�@TPA� �Q�TXa�t\j�@E�L�BM250`0/D8���$78�monf�195d SD95\F�UEC 0OP� UFQR@ ��;!C@ \�@�;!O�0pt"VIP��@#� I�@0�!CsSX� �#WEB �#HTT \st2B24 �#CG�Q#{IG�Qtopm�PgPGS!��PRC�@FSH7���w!6( B�8��![�R RBB�- Ci�B01ro�gw!#IF#"09�8-!!` �@�A64:�(AaNVD�!Ld�1h 6a68( c�`�d SR7c!te.p� 0kaч@�bc`� CLI$0?�sb$c9G MS�"5a�` w- A� STY�@wal �@CTO �CJNN0J98�ORS�0G��b��g J�`OL�1A{bn: SENDu�to�!L�Q���@*r�#SLM� 8�"F�VR� MCHN0C9SW!SPBVP�і PL� ds �qV$0�cCCG $p�aKCR�0
Np�QB� �87.f�QK� j�70*`�p�0'3CSnqToo�CTQL���qTB�P�N���@n;pqC�@�Q#�� �p,#�p ��. �%�$07#%� `8D#TmC� QSQ"TE� �[#m� �tTE� g0t"m�P�TTF�Q[�8���@�#CTG�Q�"8���@�#CTH `�T�TI�@#CT'Qe;qs�PCTM�@SC��$0gS��0bod�yqP�@  �<�� �1� 1d��q�aus�a9�H�P[�qW `@06; �GF `8�V@VP2�@ 623R i��@jH?�g� `n�g�B `�" g�D `��g�F�X mna"PVPIH��+ G V�!#V	`o  23�RVK�@,Np�@CV�Q31��934.�vo =R�erne땗�H���i��r���h���A����37� ��"�\srv����b�3b^�- Sr�B"0x���A�J935땼�B�5 (S�O@���g �1�1�R|�j93땷b���EN�5�� aw�m�SK� Lib������� �����	 �"|��h�h�#��b�wm�sk�nE����ql���pyE�  ���!�02�t F�uïբ6ۯm��u�ji-�I&���8 k��8!�Ń�땼P���2�2�2�Mai'�on��_�/r�;pڦh;�;�G��_r؈��!��4\ֶOR�C��+�5�� "T�¦TP��hQ�65�2�1��4���<�xkP�����ߦ�t�P���QrֶSB�� ch_����)�t!0�B�"
̿ h�h땇�;��� c������������x>�Rp� \toֶ�3���cl�W��2 p�"���������� F����b� Qt�a$�϶0t��ܐFsȒ��76�p�t	� A9d���582��ob��|*{�\a��FMQ ���A��migֶ�I�or��wI�j�rfm���Fc���@1�E�YE~� w���R����4�K2Х70r.�E�ld,�lC�� 1PTP]����.�"AD.�F��&3 k���ask���ȍ`4���۳d�ֶے��ER~�7 R�ƫ/�T�?)�e�rv�G?Y?k?}?8�?�?ӹapa��	�d����r�4�M��t�e����79!J�dd/���G�p�ac� T��<6�b�/� QO�&�$vc>�,@Vg��"��eYW��5/�c BJ�h���R5:�d���0�@��I_��raj��e��hQe}�$`��5(Xa�@Ƈ�et榻�1Otd�j��,�_h�\	UI�/k�jo�FO��`�^���F��r��qW6�5q���K �'6ڦu7s W'�b,'��t'?��n��MFR�ֈ;]�lf�ǯ�fr>֛�w�p�/�,@��_U[ǀ�мn�x '_i�{�����O���p`J���[@�o�in7�L�O�9�\^ � R����+mi2״h �j��҇;- f�nt >��MA H�I  H5529ķ (Cߑ21��l?eR78�c��ߒ0AcaJ�614���0A�TUP�����54]5�t-fl�6yE�=�VCAM�tFL?XCRId����o�UIFULX ��28��mo�NREu'��63��WQ���SCH��Cn�DOsCV�gϠCSU1��cxr�0$�;�EIOC%tx\�c��54�oQ��9�T�;�ESET�TeCmo?�S�/��7S��{�MASK��70��PRXY�T�`���7��`�OߐOCO
e�\?�3�ô`>��!0{�?��|�-��oon G?�39!'�ߑõ H82�LCHd��@I�OPLG�tCGM�?�0��GЎ�MHC�R�Go�S�/1_�C�S4�cgm��50�T��?�5$�[���M'DSWMf.�D������OP��X/2L_�PR��K�����{����883n�CM^��0iA,��0����`~�5#�\h88@�+�?�D���.?�*��4��0D�3��o��S4����9��,i�FRDd�/2�E/��MCN5�H�93�K�SNBAv�U"R��HLB�ɃSM�՛ñ�T���Jc52�SaߐTC4��\�TTMIL�e��P���A|�TPyA���TPTX�ŝ5��TEL�ԫ�0䴈P��8�˳���fK�95����95��w888��UECd�wrt �UFRd��__�Cd�2e-�VsCO4��VIP�;��I�TAX~�C�SX�����WEB84����HTT4�kaz��2T�2M/So�yG#��QIG��< .�IPGS=t\rxO�RC��aߐ7�/a��6D�s@>�R7#��!��Oq�� ���P��Ҷ;�A���K�\��$�0 "��4�����NVD4���#�A�dap��8D���68����R7���P��D0��a��o�bܠn. CLI��l\-C���CMS�'���4�d "ްSTY��[�CTOT�tl枱NN����ORSp4�;�1 ��ltiΰOLS�( E���0�T���L��6�@����9@ ��LM4�HV� o�VR���C�S��shc>�PB�V4䫁/�PL�
A�PV��ust>�CcCG4��0nCR�/4 H5��B��z�K�H573����?����\cms��#�st.~TB����! ��7�C�ԓ�?"�awshD?"��I0?"��3��TCd�K�A 4�\sl"EĤpP��� 4�C[П"Ԥ8c��"4�\(��CTF��c���"���CTG�7e3m#G�THd��h� �I��K�CTvC�59m�CTM��5M����Q0��re\g�P���12���04�����%Sv��13MCTWd��9[@_�GFd�SE]�P2d�t+��2�ո� �2d�ell��P%Bd�I���1Dd��a��1F��tap V3PId���CV�!�Vq��UA��CVK��ۣCV#�cor�eL���H"�Hpp!�HK"�Hatc�JH�H�4�I� �IL0H�I�2�H��H+2�IL�Y4=�H���I�e\a�I�2 Z93��I{�H�@NZ+��H �1��K48�Z<A�Ht�{�Il �Z;"�O�Fs \!�Hk"�H{"@o�F[�BPZo�Z���J��Tok �РH��H\��Il�hZ��Z2=[ng-[gToo�I�p�j(��njrobt_�Xbct.�JL� iur�o��I��i�!��F��POz�ling�j��y���Y"r^zۢ�I�p��Geat^j�]��Z��_je�����_��lkҠHm,��H|���Z��A�I  ��_�  ���Gvhm�J{�svnj���H�49\�J�@L�Ij�749{P�Zt\ajNj�@_"g.pj�mcal�0�fu�J��^zhm-��_bg(���o�\ͫ �1�H�! j��;����MT; "�(Cu�zkL��bgft�JlpX����GCT"���Gfyc]�˝26\fߟ�926�l\� Ί�u�>m��;�Mu1l?�Q��7\^�K����7-[˝���_�6�1Nj48.� H�- �H�@R_�L^zi�Pe��K�Я�F8\�}�}�����Ћ� � yRk,�ticMoj+@OoQxs-@�"�3�gCS j+}LB-[�5 HNj+� co�~�L��z��f�k˝lb�jll����-˂��k/�.���LЎ�kwipJ/�on,�Jt\A��8�SK"��� ��uto�o aB������kwm�1 �o��Htp�ʜ �n}��ex-�˝��x����a^jlL�je$�식i��a��/����rej�1��o�Vor�zR����e T�Z[��[GlclN��߭�SOz�̌GZD��to8�{+B�H643N�`�cSG/o��sg�a�Utui��;`�J���`�;�ndm�ndiN�{/�/�/�/�/ �/�/�/??/?A?�?���riΪ! -Kj7950/�n �zk]�895n/�O�t �Z��wsg�K,�>���iag� SG8J�Ю�ogu����KO]Ltw>_@	J6�4�1�s�{F O�>ګcdݛ��`3d_��r-��N74�uy-�3��RINnzlly��(m^���Lܬ��sgc�zI"� #?
+�oߡ\tw/��0.�@�"���(f�_�[y�Kmm�K}�dct^�t]�+�
{PRZWCHK
�k,�;;`y<p��l�K���LN*R852j �@_jR ����tiN�g WJh�ecN�L�F����w�lZ|*�da9t�ʛ�greN���o  S�TD�r7L�ANG�Aoc�e��`��Q�7��R�870�{��8 {(P�ogge�p��!�58\㕏PATTs�� �t9\��c "B�@�V��1�patd���O���������({q㕔�5�a�p[��m�\㕻�7�\aAw��@�a��p6�𫯽�ϯ�gmon���d��0�B�m�@;A��\ ö��K�I��MHCR�51 	H����g\o��@��=R]� H54ۿm�<@E���;!�����Gomm�;a��R�"|�N㕬0F�C��W�P�)Ai6�� Fƫ�\{��itx�#{ ���iaio����D�e6�eve����7C2 R�@RƜPg��7adl��nt��K�RBT�t�OPTN`772'�CTK"'�g�(�x���)� "AZ'�p;q'�q'�tzn&�{ E'�Ama��-� Mu��ncInDPN����<���872��|�d��(��������#���masy��y "M��o��䃲��#et����\p1������\ ��f���lZ ����lp���9���`p��+ V��ail��@?��䇢�䓢��zd�x<�k`��73.f���irdg��- i���e\ ����� S]0j�021"�1W ��(�`�4�� (i6��e,"� "���+���core_�I���l`F��AY��AB��@����H������ABIC��Par;�M�ai�������<� c\�ITX�>���  ����w1��g Jcwlib��Shi�W�4�� t994\�VSSF��� t�t\j9�f "�O�w� t��$%ini�/��pٰ t�p5G�&,� t\vsR&�x�L�%w� tamcylS/+ref.�%$#� tj��%m�� t�[A�&4\z�/�,z�_v�%A�%�a�%_�ol6��l% �%end�/<c?.?@?�R5o[?m>�6�/�dsshf�/+trt�?�<OAE�'F  !`�G��$%��5vi�6<���6 J92�F3���%25 (�%�@e�&�P�%k�4O dn�wzF��T�&`�XEp�n�&g��? nw\�n�?�,nd�V��N�;XnF j���%se�V I/
&�q&Ѹ�U��5r w�%/aF� �F�_�rclR&�0\pw/Y�90�E�o`/"5Of "U<//A+dprm�%g��%�Xrsu/kmS�T_! L`�6/OŔpM�LO��j��nO1|h�ODn�on�|YCwrp�R/�l���E<�Pe\gya��Krgas�o��k��f�v��4x1tf�?m$ra�o�l�a0�omk�_�Tam�N6+�4�`'9K0.Av�Wې�%�@�Ft���XE sV��ДJ7{37�%|*�%�,P��hB "+��Kw�cfF& I����9�98�vtomzFut vV�_	o;�YC����:8\F&�Y/� t0��f��deb^V ��$�0zFؠ"�䠙g���<9\�&��9��Wr}  �su"�s�t�G��X �f� U (�fagn�F PzFlϜ�Via�TX����vd��w��g��HnzF- O�W CH� �$723�F���E(A�ÿտ2蚽Wc�6�WsvF& S�W�J�R6��_�RVo `RV���ӊ��vt��M\etF�XoN�o��Fr��x���+�1T��F?teR� J5�8�O  34	Wg�le,�%,�j�Dq\at"��zFwIta1FlUTA�VϜ�gw��Mad�W�Oa���6d M��e�FT��o90 H�%NT��R69������i;r\ʆMIR��ӊenʆv���F|�3�N�ITCP��Ta0�p���(MM7G�eT^�o \tpʆI��NYBbusJ׈�m� �I�@zFȀ��F������/��W�'g, 0��4`R_(!sw�&s_�YC67\JF��Tf1_����Dfw��W�Ι4achg��a96�_��� _���_r�V�% 9�9YA�e��$�FEAT_ADD ?	������  	 �$YA//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ��߿������DEM�O N�   ��*� �2�_� V�h���������� ����%��.�[�R�d� ���������������� !*WN`�� ������ &SJ\���� ����//"/O/ F/X/�/|/�/�/�/�/ �/�/???K?B?T? �?x?�?�?�?�?�?�? OOOGO>OPO}OtO �O�O�O�O�O�O__ _C_:_L_y_p_�_�_ �_�_�_�_	o oo?o 6oHouolo~o�o�o�o �o�o�o;2D qhz����� ��
�7�.�@�m�d� v�������ƏЏ��� �3�*�<�i�`�r��� ����̟����/� &�8�e�\�n������� ��ȯ�����+�"�4� a�X�j���������Ŀ ����'��0�]�T� fϓϊϜ϶������� ��#��,�Y�P�bߏ� �ߘ߲߼�������� �(�U�L�^���� �����������$� Q�H�Z���~������� ������ MD V�z����� �
I@R v������/ //E/</N/{/r/�/ �/�/�/�/�/??? A?8?J?w?n?�?�?�? �?�?�?O�?O=O4O FOsOjO|O�O�O�O�O �O_�O_9_0_B_o_ f_x_�_�_�_�_�_�_ �_o5o,o>okoboto �o�o�o�o�o�o�o 1(:g^p�� ����� �-�$� 6�c�Z�l��������� Ə����)� �2�_� V�h���������� ���%��.�[�R�d� ~������������� !��*�W�N�`�z��� �������޿��� &�S�J�\�vπϭϤ� ����������"�O� F�X�r�|ߩߠ߲��� �������K�B�T� n�x���������� ���G�>�P�j�t� ������������ C:Lfp�� ����	 ? 6Hbl���� ��/�/;/2/D/ ^/h/�/�/�/�/�/�/ ?�/
?7?.?@?Z?d? �?�?�?�?�?�?�?�? O3O*O<OVO`O�O�O �O�O�O�O�O�O_/_ &_8_R_\_�_�_�_�_ �_�_�_�_�_+o"o4o NoXo�o|o�o�o�o�o �o�o�o'0JT �x������ �#��,�F�P�}�t� ������������� �(�B�L�y�p����� �����ܟ���$� >�H�u�l�~������� �د��� �:�D� q�h�z�������ݿԿ ��
��6�@�m�d� vϣϚϬ�������� ��2�<�i�`�rߟ� �ߨ���������� .�8�e�\�n���� ����������*�4� a�X�j����������� ����&0]T f������� �",YPb� �������/ /(/U/L/^/�/�/�/ �/�/�/�/�/ ??$? Q?H?Z?�?~?�?�?�? �?�?�?�?O OMODO VO�OzO�O�O�O�O�O �O�O__I_@_R__ v_�_�_�_�_�_�_m  h$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲�����������   ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ��������
��	�,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_�oi�$FEAT�_DEMOIN [ d�D`�`},dINDEX9k�Ha�,`ILEC�OMP O�;��zaGb'e�p`SETUP2 �Pze�b��  N �amc_A�P2BCK 1Q~zi  �)hD�o�k%�o`}` Ae�om�o�  ��V�z�!�� E��i�{�
���.�Ï Տd��������*�S� �w������<�џ`� �����+���O�a�� �����8���߯n�� ��'�9�ȯ]�쯁��� "���F�ۿ�|�Ϡ� 5�ĿB�k�����ϳ� ��T���x��߮�C� ��g�y�ߝ�,���P� ���߆���?�Q��� u����:���^��� ���)���M���Z��� ���6�����l��� %7��[���  �D�h��i�`�P�o 2�`*�.VR`� *�c�����JP�C��� FR6�:�.�4/�T X`X/j/�U/�,;`%/<�/�*.FM�/"�	��/<�/<?�+STMG?q?��D]?�=+?�?�+H�?��?�7�?�?�?EO�*GIFOOyO�5eO"O4O�O�*JPG�O�O�5`�O�O�OM_�JSW_Ā_� Sn_+_%
�JavaScri3pt�_�OCS�_o��6�_�_ %Ca�scading �Style Sh�eets0o� 
A�RGNAME.D)T_o��0\so1oГQ�d�o`o�`DISP*�o�o�0�o7��e)q8�o
TPEINS.XMLg�:\{9�aCu�stom Too�lbar��iPA?SSWORD.�?FRS:\��� %Passw�ord Config@��������� ��r�����=�̏ a�s����&���J�\� 񟀟����K�ڟo� ������4�ɯX���� ��#���G�֯�}�� ��0���׿f������ 1���U��yϋ�ϯ� >���b�t�	ߘ�-߼� &�c��χ�߽߫�L� ��p����;���_� �� ��$��H���� ~����7�I���m��� ����2���V���z��� !��E��>{
� .��d��/ �S�w�< �`�/�+/�O/ a/��//�/�/J/�/ n/?�/�/9?�/]?�/ V?�?"?�?F?�?�?|? O�?5OGO�?kO�?�O O0O�OTO�OxO�O_ �OC_�Og_y__�_,_ �_�_b_�_�_o�_�_ Qo�_uoono�o:o�o ^o�o�o)�oM_ �o��6H�l ���7��[��� �� ���D�ُ�z�� ��3�ԏi������ ��ßR��v����� A�Пe�w����*����N�`���֦�$FI�LE_DGBCK� 1Q������ (� �)
SUMM?ARY.DG����OMD:3�s����Diag Su�mmaryt���
CONSLOGi��L�^�������Co�nsole lo�g����	TPACCN�R�%:�wς��TP Acco�untinρ��FR6:IPKD?MP.ZIP�ϯ��
���σ���Exc?eption ߱��_�MEMCHEC�Km�Կb����M�emory Da�ta��֦LN�=)n�RIPE�\߸n���%�� �Packet L�Ϻ��$SA���S�TAT�����ߋ�� %�Sta�tus��<�	FTAP����r������mment TB�D��� =�)ETHERNEU����B�S�����Et�hern(��fi�gura߇���DCSVRF���������� verify all�٣M(��DIFF����/diff�PB���CHGD1�x�� �FQ&���	2��� 5�YGD3p���'/ ��N/�UPDAT�ES.m S/��FORS:\k/�-���Updates �List�/��PS�RBWLD.CM��/���"�/�/�P�S_ROBOWEyL1���:GIG����?/�?��Gig�E ��nosti�c*�ܢN�>�)}�1HADOW�?��?�?5O��Sha�dow Chan�ge��٤&8+�2NOTI��O"O��O��Notif�ic��\O٥O�A��_��2_կ?_h_ ���__�_�_Q_�_u_ 
oo�_@o�_dovoo �o)o�oMo�o�o�o �o<N�or�� 7�[���&�� J��W������3�ȏ ڏi�����"�4�ÏX� �|������A�֟e� ����0���T�f��� �������O��s�� ���>�ͯb��o��� '���K��򿁿ϥ� :�L�ۿp����Ϧ�5� ��Y���}���$߳�H� ��l�~�ߢ�1����� g��ߋ� �2���V��� z�	���?���c��� 
���.���R�d�����������$FIL�E_� PR� �����������MDONL�Y 1Q����� 
 �)�@_�VDAEXTP.�ZZZ��p�G�L�6%NO Ba�ck file <!��U3�M�� 7����G�&� J\����E �i�/�4/�X/ �e/�//�/A/�/�/ w/?�/0?B?�/f?�/ �?�?+?�?O?�?s?�? O�?>O�?bOtOO�O 'O�O�O]O�O�O_(_~��VISBCK��|��*.VD)_|s_�@FR:\BP�ION\DATA�\^_R�@Vision VDt �_�O�_�__o_Ao �_Rowoo�o*o�o�o `o�o�o�o�oO�o s�@�8�\� ��'��K�]���� ���4�F�ۏj���� ̏5�ďY��j���� ��B�ן�x����1����ҟg���MR2_�GRP 1R����C4  B�O�	 
������/E�� ֯�r����OHcEP]���O��#M��^
�KA���?��&�r���:6:�N�R�9-�<Z��A�  v����BH��C`}dC���N��B�{���r���пὫ�@UUT��U�����/Ϫ�>��>c���>rа=����>i�=����>����:���:��:�/:6)�:��~ϗ�2ϔ��ϸ�������z�_CFG� S��T � �a�s߅�0[NO {��
F0��� ��/\RM_CHKTYP  ���O����������O=M��_MIN��L�g�����X���SSB7�T�� ��5�L�,�U��g���TP_DEF'_OW��L�����IRCOM�Ѝ���$GENOVRD�_DO��	��T[HR�� d��d��o_ENB�� ��/RAVC��U�UQ �Υm�X��|��������� �� �OU��[���O����⾥8��:���
,.  C�x �h�������B�ϡ������n�!�SMT'�\�.���+�w�$HO�STC7�1]K[��Y��� MC�L��MI��  27.0�1�  e}�� � /*�1/C/U/g/��!/#	anonymous�/�/�/��/�/? L��8 ;{}/j?��?�?�? �?�?/�?OO0OS? �?�/xO�O�O�O�O? UO+?=?_QOs?1_b_ t_�_�_�?�_�_�_�_ o'_]OoOLo^opo�o �o�O�O�O_o G_ $6HZl�_�� ����o1o� �2� D�V�h��o�o�o��� ԏ��
��.�uR� d�v�������?��� ����*�q������� ����ݏ��̯ޯ�� I�&�8�J�\�n���ǟ ٟ��ȿڿ���E�W� i�F�}�jϱ��Ϡϲ� �ϋ�������0�S� Tߛ�xߊߜ߮���� �+�=�?��s�P�b� t����ϼ������� �'�]�o�L�^�p������/ENT 1=^�� P!���  ������ *��Nr5~Y ������8 �\1�U�y �����4/�X/ /|/?/�/c/�/�/�/ �/�/?�/B??N?)? w?�?_?�?�?�?�?O �?,O�?ObO%O�OIO��OmJQUICCA0�O�O�O_�D1_�O�OV_�D2W_3_E_��_!ROUTE�R�_�_�_�_!P�CJOG�_�_!�192.168�.0.10�O�CC�AMPRTGo#o!�7e1@`noUfRT��_ro�o�o��NAM�E !��!R�OBO`o�oS_C�FG 1]�� ��Aut�o-starte�d��FTP�� ~q���F���� ����9�K�]�o�� ��&���ɏۏ����� Wi{X����o��� ��ğ֟������0� B�e��x��������� ү�������Q�>��� b�t�������q�ο� ���9���L�^�p� �ϔϦ�������%� �Y�6�H�Z�l�3ϐ� �ߴ�������}��� � 2�D�V�h�������� �������
��.�@� �d�v���������Q� ����*<��� ���������� ���8J\n� �%�����E Wi{}O/��/�/ �/�/�/��/??0? B?e/�/x?�?�?�?�? �?/+/=/�?Q?>O�/ bOtO�O�O�Oq?�O�O �O_'O(_�OL_^_p_��_�_(�`_ERR� _z�_�VPDUSIZ  9P�^S@��T>�UW�RD ?EuA��  guest3V$o6oHoZo�lo~o�dSCD_GROUP 3`E|� Iq?YM ��nCON�nTAS��nL��nAXP�n_�E�o9P�n�RTT�P_AUTH 1�a�[ <!i?Pendan�g�~�@}9PJ�!KAREL:*���}�KC����p�VISION SCET�`E��I�!\� J�t��s�����������Ώ��-���dtCT_RL b�]~��9Q
@<FF�F9E39�DF�RS:DEFAU�LT��FAN�UC Web Server����bv odL��'�9�K�]��o��TWR_�`FI�G c�e��R���QIDL_�CPU_PC�9QB�@� BH�ǥMINҬ�a�GNR_IO�Q�R9P��XɠNPT_SI�M_DO�!�S�TAL_SCRN�� �y�+�TPM?ODNTOLY�!���RTY8��&�9�.hpENBY��cƣOLNK 1d�[�`�����1�C�|U�ͲMASTE����&�OSLAV�E e�_˴jqO�_CFGsϦ�UO�D��Ϩ�CYCLE��Ϧļ�_ASG s1f���Q
 W� 9�K�]�o߁ߓߥ߷� ���������#�_��GNUM�S�b�U
���IPCH��j�O_RTRY_CN���Z��U�_UPD�S���U �����g�θ`��`ɠP�_MEMBERSg 2h��` $�e��>��HyɠS�DT_ISOLC�  ���r�\J_23_DS��q�~��OBPROC��n%�JOG�d1i���89Pd8G�?�.���.�?�?�?OQNs��V ����3W~�����������POS�RE��$�KANJ�I_m�K�i�pMON j�k~�9Ry����//�^$�r��k����9%Th��p_L�I�l�k�EYLOGGINʴ��`����U��$LANGUAGgE �����Y �!�QLG��lq��9R��9Px�p� � ��砬9P'�03X�k���M�C:\RSCH\�00\��� N_D?ISP m��DpAMK�SLOCw��آDz ��A�#O�GBOOK n���9P~��1�1�0X�9O%O7OIO[O�mN�Mɱ���I��	��5Ib�5�O�O�5��2_BUFF 1-oؽ�O2A5!_ �2��=_?7Y_k_�_�_ �_�_�_�_o�_o:o 1oCoUogo�o�o�o�o�e4��DCS q>�= =��͏L�O�-�1CUg���bI�O 1r� ��s20���� ����1�A�S�e� y���������я���@	��+�=�Q�|uE�TMl�d����Ο �����(�:�L�^� p���������ʯܯ�p ���7�SEV��u={�TYPl����z�����!�PRS����/S��FL 1s�}����$��6�H�Z�l�~ϯ�TP� l�i��=NGN�AM��A5�"e4UP�Sm0GI��\!�����_LOAD��G� %u:%PL�ACi�2�3�MAXUALRMI�c�W�T���_PR���h�3�R�Cp0t�9��M���3Eݗ���P �2u�� �1V	Zi�00���� ��1��.�g�xU� ����������� ��8�J�-�n�Y���u� ����������" F1jM_��� ����	B% 7xc����� ��/�/P/;/t/ _/�/�/�/�/�/�/�/ �/(??L?7?p?�?e? �?�?�?�?�? O�?$O OHOZO=O~OiO�OK��D_LDXDIS�A����zsMEMO�_AP��E ?��
 b��I�O _"_4_F_X_j_|_RпISC 1v�� ��O�_ ���_�_��Ooo@o�_C_M?STR w:�_e�SCD 1x�M� 4o�o0o�o�o�o�o P;t_�� �������:� %�^�I���m������ ܏Ǐ ��$��4�Z� E�~�i�����Ɵ��� ՟� ��D�/�h�S� ��w���¯���ѯ
� ��.��R�=�O���s� ����п����߿�*� �N�9�r�]ϖρϺ��PoMKCFG �ynm����LTAR�M_��z������и���6�>�s�MEgTPU�ӫІ�vi�ND��ADCOLxXի�c�CMNTy�s l�g` {nn���-�&�����l�PO�SCF����PR�PM����STw�1�|�[ 4@�P<#�
g��g�w�� c���������� ���G�)�;�}�_�q������������l�SI�NG_CHK  �|�$MODAQ��}�σW��#DE�V 	�Z	M�C:WHSIZE��M�P�#TASK� %�Z%$12�3456789 ���!TRIG +1~�]l�U%�\!��S
K.�S�YP�69"EM_�INF 1�� `)�AT&FV0E0�X�)�E0V�1&A3&B1&�D2&S0&C1�S0=�)ATZ�#/
$H'/O/�Cw/(A/�/b/�/�/�/? �&?�� �/�?3/�?�/�?�? �/�?�?"O4OOXO? ?�OA?S?e?�O�?�? _CO0_�O�?f_!_�_ q_�_�_sO�_�O�O�O �O>o�Obo�_so�oK_ �owo�o�o�o�_�_ L�_o#o��Yo� ���o$��H�/� l�~�1��Ugy� ��� �2�i�V�	�z��5�������ԟPNIwTOR��G ?k�   	EX�EC1���2�3��4�5�� �7*�8�9����� �����(���4���@� ��L���X���d���p����|���2��2��2���2��2��2Ũ2�Ѩ2ݨ2�2��3ʉ�3��3(�#R_�GRP_SV 1݀� (�ſ1�x�>Ka����?|���R��_Ds����PL_NAME !����!Def�ault Per�sonality� (from FwD) ��RR2��� 1�L6(L�?����	l d��nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲�����B2]���*�<�N�`� r����<���� ������,�>�P�b��t�����BJ � �\  ��  �����  A�  B��UT��� 
����~���  �������B��p��� � CH CH P �Ez  E�� E�` E��;%�Z��*� �  E���F�@&�U�T Ai�  dx�H�x�	$�Hxd�dڭ� }`(d��8�(xx$$ y Xtd D (DDdpWwX� �	X�vXHX����/y�y (�� !��  7%E	��Em�Xw�$%XH$%P��  �/�/�/�/�/�/??�+?=?O?a?s=F��r?�?�?�?�6��E�2ExB�2
�������?Kزd��'O9NO\OjG��0��|M��ն'4� � W%8�O�O�N �0�G��O�JA  A��C�����_�OC_9W�
  � TB�LY��
��_�\��Q�Y=�C�و�V�`HR0� ʒ_P( @7%?���a�Q?ذaر@��6�&س��2n;��	lb	  ����p�X��U�M`��X � � ��, �rb��K��l,K���K���2KI+�KG�0�K �U�L�2o�E	O�n��@6�@ t�@�X@I��b`�o��C�N����
���}v��#���` q�m�|�kQ?�
=ô��  �Hq�o`!b���9�  ���a� �� ���ذa�s�G��}2�m��o�q��v�O���E	'� �� 0�I� ��  � Q�J:��ÈT�È=��9�l���@|��� }~�Q����R������N8���  '���ap?��P�b!p�b){�B���?�CIpB  X���ذ��C�A�a�/ � {��	�o�Q�IB P��8�����P��ԕرD �O���O���A�,���Š
�`l�1�	 �٠p��� p` rl`:�4  �t�?�ff{O��įV� �P�����a�,!�/�?Y)R�a4�	(ذ]�Pf����a\c�\dƃ?333-d����;�x5;���0;�i;�d�u;�t�<!� +}�oݯ��b�Sb��P?fff?��?�&��T@��A�#$�@�o[ ,ž�x�	�&f6�ed� g���Hd㯸ϣ��� �� ���$��H�Z�E�~߾�&eF��mߺ� i���U���y���2���E�0����y�d� ������������ �?�*�܏r�8�.o�� �����T�); ڿPb������0��P��A��T C�=�ϵ��Y}��2��������C��W�C�>= �` Ca���B����(!�`�<����bC@_;C�9�BA��Q�>V{�������Y���uü��
/��S��Q��hQ��A�B=ן
?h�Ä/iP���W��È�K�B/
=�࿣��Ɗ=�K��=�J6XK��r#H�Y
H}��A�1��L�jL�K���H:���HK��/0	b�L �2J���8H��H+UZBu�a?�/ ^?�?�?�?�?�?�?O �?O9O$O]OHO�OlO �O�O�O�O�O�O�O#_ _G_2_k_V_{_�_�_ �_�_�_�_o�_1oo .ogoRo�ovo�o�o�o �o�o	�o-Q< u`������ ���;�&�K�q�\������Gϭ���� �C�aɏ Ĉ���CVF������+b����Kc�f�� 
E�����T�ٟ�(��g_�h۟�������N��������3lC�(�:�H����T�f��t�.�3��}����k����q'�3�JJ�����گ���4��"�]P̲Pf��� ����⟛�ſ���Ի�����/��?�{x?�N�u�  fUh� *ϳϞ������Ϣ�t�0.��R�@��X�bߘ�߆ߨ�)Z�ߺ� ? ( 5�	�߀����B�0�f�t�  2 E%p"�E[@��N�"BXC��%@ߏ��%������)�;��������������%n�n�%"��%��Xc
 ��!3EW i{��������b*[��P�I��v�$MSK�CFMAP  ���� �^�����pDONR�EL  X��[��DEXCFE�NB�
Y�F�NC��JOGO/VLIM�d��]dDKEY��=%_PAN�"\"DRUN���>#SFSPDTY�w����SIGN|��T1MOT���D_CE_G�RP 1���[\���/��?&?�� ?Q??u?,?j?�?b? �?�?�?O�?)O;O�? _OO�O�OLO�OpO�O �O�O_%__I_ _m_�_f_�_O�DQZ_�EDIT�$UT�COM_CFG 1�Q�_o"o}
�Q_ARC_��X��T_MN_gMOD���$�UAP_CPLFo��NOCHECK� ?Q  W����o�o�o�o '9K]o������vNO_WA�IT_L�'�W� NMT�Q�Q���o_ERR�!2�Q��� �_t��������*��Ώ�d``O�I��P�x b��_���8�?���4�����B�PA�RAMJ��Q����	�����s�� �=��345678901��� ���?� Q�-�]�����u���ϯ���������7�~ODRDSPEc��&�OFFSET�_CAR�PKom�D�ISz�K�PEN_FILE���!$a�V�<`OPTION_�IO
/=!аM_P�RG %Q%$�*	�ά�WORK� ��'� C��Kƪ�P����Ɋ��f�(�f�	 a���f�5���M��RG_DSBL  Q�����L�RIENTTO* ��C���Z��M��UT_SIM_D�طX+M�VQ�LCT �%��R_�x$aQ�'�_PEXh`ܜ�b�RAThg d�b�r�UP )�5� � �����X������$��2�#��L6(L?}��	l d'� O�a�s������� ������'�9�K�]�@o���������H�2>� ����/ASew�N�<����� ��1CUg�yH���P��� �  �� � �U�A�  B���PB�����H��  ����U�B�p�������N�P E�z  E�� E_�` E��;(�����Z�/�~��  E��''l���@#���T�AJ(��E!Y! a!)!m!Y!u)%)!Y!(E!�%E!ڎ$�^$A! �	!E!a!�%%	-Y! Y%�-58�Z 99HU%E!�D!	$D%% E!Q481X291�%�)95 �/W#95)%91m5a!�5)/Z7��Z (�8�1a�<a1 EE	�(�Em�494X6E9=8)%E15�� |O�O �O�O�O�O�O�O__80_B_T]F�S_y_ �_�_�Vh�����_�[��%�on�_=o�Kg�]�]&�'4 � W%po�oX� ���g�o�j�A�A��c������o�o$w���tB�(~�`��r�|B�� q�y�$�O���1�'k�'ۆ�3�`��0���P�( @ED�D��q?�Q�C�Z7}��o  �;�	lD�	u� ����p�X�[�2���X � � ��,i�X��`H���9H�H����H`�H^yH�R�l���_h�����`C#�B�� C4ӄ����c��9���
=���� ������c�Bz��Βa�m�另b��s�� �q���g䟒����Ǒ�ٖ�o���e	'� � ��I� �  ��q<�=���89�K���@a�g� b���������唠�䮟�N��  '۰��Ɓ"�B�Ղ���т6��� �  O��C�a��	m�~��p=�Bp��Н� ���px����D��o�޿�o��&��o��5�Ю`Q��	� ٠U�f� �U� Q�:���#�>���?�ff\o����;� �p����"��8� ��?Y
r�$�q=�(� B�PK�f����A�A���?333���m�;�x5;���0;�i;��du;�t�<�!��y������t����r�p?fff?�x�?&���@���A#	�@�o[�	]����� �uI��wh���-��ϝ� ���������	���-� ?�*�c�u�L��������4�V�X����EjPf��^I�m ���� �$ ��W������ �9��/ /��5/ G/�z/e/�/�/�/�/��`�A��$�t�/ �C�/"?�(d��>�?��Pn?�/�?}?�m�(��W�?C�@�` CT��?�j4�j0i1A@I��!���bC@_;�C9�BA�Q�>V`.�È����Y��uü��
��?�3��Q��h�Q�A�B=?�
?h��iOJp���W�����K�B/
=����Ɗ=�=�K�=�J6X�K�r#H�Y
�H}��A�1��=L�jL�K���H:���HK��O�@	�bL �2J���8H��H+?UZBu�?F_ �OC_|_g_�_�_�_�_ �_�_�_o	oBo-ofo Qo�ouo�o�o�o�o�o �o,P;`� q������� ��L�7�p�[���� ����ȏ�ُ���6� !�Z�E�~�i�{����� ؟ß��� ��0�V�8A�z�e�Gϭ����� C�a�/�� �爓�ЯׯCVF������üKG�j����KH�K�� 
AEp�s�9���90(91ϳ_�h��y���<�i��N����T�3lC���-���9�Kϰt��.3��}e�w�k����q'�3�JJ�͑��Ͽ�����(��B5P��PK�Zgt�ǿ�ߪߕ�������������$��{$�3�Z�  fU M���������`Y��7�%��=�0G�}�k���)Z����  ( 5��  ������'KY�  2 E%pnIFE[@tN�IF�B�!�!� C��0� T�@į����*H3��Tf�x��T�T�"94��T�D=4H;
 �//*/</ N/`/r/�/�/�/�/�/��/�/GJ@2��5�I��v�$PAR�AM_MENU �?����  DE�FPULS��	�WAITTMOU�TT;RCVg? �SHELL_�WRK.$CUR�_STYL��Γ<OPT��?PT�B�?�2C�?R_DECSN_0<�L	O O-OVOQOcOuO�O�O �O�O�O�O�O_._)1�SSREL_ID�  ��Y�=UU�SE_PROG �%8:%*_�_>SC�CRk0ORY@3�W_HOST !8:#!�T�_�ZT\Ю_� c�_�Qc<o�[_�TIMEi2OV�U~)0GDEBUGMP�8;>SGINP_F�LMS`�gn�hTR\�o�gPGA�` �l�C�kCH�o�hTWYPE5<A)_ #_Y�}���� �����1�Z�U� g�y����������� ��	�2�-�?�Q�z�u� ������ϟ�
��eWORD ?	8;
 	PR�`�U�MAI@��3SU�1E�TE#`U���	�4R�COL�S�n���vTRACECTL 1��ŻB1 W 6 7�W d�ެ��_DT Q�����РD � *������W.��.��.���`.��"��	��
���
2�:�B�B����"���;���3�:�B� J��+�=�O�a�s��� ������Ϳ߿A�S�a� �[ÑĠϲ����� 9�������	��-�?� ̨ߺ�����P�b�L� ~ߐؓ���)�;�� '�Y�k�}�oρϛ�� ����������+�=� O�a�s����������� ����'9K] o�0\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz�uX��� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��ߚ���� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p����� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�?��?�?�?�?�?OA��$PGTRACE�LEN  A � ���@�$F_UP _����SA[@�?AT@$A_CFoG �SE=C*AT@��D�D�O�G6@�OhBDEFS_PD �sLA�6@�$@H_CONFIG �SE�;C @@d�T�3B AQP��D�A1Q@�$@I�Nk@TRL �dsM�A8�EFQPE�E;�W�SA�D\Q�ILIDlC�sM�	�TGRP 1��Yb@lAC% � ��l�AA��;H�N��R����A!PD	� a3C	\T�Ai)i�QP� 	 p�O4VGgCo ´|c^oGkB`�a�opo�o�o�o�o�b"�B�z�o7I~3 �<}�<�o N�J����� f�)��9�_�J�`z����@
t���d� ŏ�֏���3��W� B�{�f�x�����՟������J)@)
V�7.10beta�1�F @����@�A&fif�Q2�CPC�`͊D�Dk`[�C��T��@ DĠ oDr� �QBH�`Y�L��PC5R Ao?�  ��CCx����b��P!P��A�����Ap�B�b!PA�1������
�?L���?333A@8��"��Fff.��bw�w:�7��A�eC�QKNOW_�M  �E{F�TSoV �Z(R �C������ʿ��ٿ��$�A!m�SM�S��[ �B�	�E���Ϗ��*�E`��2�E@�2��������� L�MR*�S�Y�T�j���A�C5����e@�Rۚ]S�T�Q1 1�SK
' 4�U��A�¨� �E��*��߽������ �J�)�;�M�_�q�� �����������F��%�7�|��Ep�2{���A�<�����PA3��������p�4��+p�5HZl~p�6����p�A7� $p�8ApSewp�MAD0F� [Fp�OVLD  SK�ϼOr��PARNUM  �/�O//T_SCH� [E
}'F!�)=C�%UPDF/X)�/|3Tp�_CMP_O��0@T@@'{E�$E_R_CHK5yH!6
?;RS�]��QG_MO�o?�5_k?~��_RES_Gz��~ݍ��?�OO�?%O O*O[ONOOrO�O�O �O�O�O�O��3���<�?_�5��(_G_L_ �3G g_�_�_�3� �_ �_�_�3� �_o	o�3 @$oCoHo�3�co�o<�o�2V 1�~կ1�e�@c?��2T?HR_INR�0�!�7³5d�fMASS6 ZwMN5s�MON_QUEUE �~�f��0��� �4N0UH1N8Ev6;�pEND�q�?��yEXE��u� B�E�p��sOPTI�O�w�;�pPROG�RAM %hz%��p�ol/�rTAS�K_I��~OCFG �h/\����DATARè��@��2�����#� 5�G��k�}��������^�ן������IN+FORé܍�wtȟ e�w���������ѯ� ����+�=�O�a�s����������Ϳ(�4���܌ �I��� K_ƒ����T��ENB� ͻ1>ƽ�I���G��2�� P�(O�ҡϳ� ������_EDIT ����ߋ�WERFL�x�cm��RGADJ �&8�AС�i�?�0t��
qLֈq���5��?�!��<@��*�%���@ؘ#ߊ��2���F�	�Hpl�G�b��>��A�d�t$�I�*X�/Z� **:c�0V�h�� �Ǟ���B������ ������������� b���L�B�T���x� ��������:����$ ,�Pb��� ����~( :h^p���� ��V/ //@/6/H/ �/l/~/�/�/�/.?�/ �/?? ?�?D?V?�? z?�?O�?�?�?�?�? rOO.O\OROdO�O�O �O�O�O�OJ_�O_4_ *_<_�_`_r_�_�_�_�"o�_�_ooo�f	 ���o�p�o�o�dJ��o�L��o#�oGY��P?REF ����p��p
L�IORI�TY����P�MP�DSP�>ߴwUT�z�4�K�ODUCT�w�8�\�OG�_TG;�|�����rTOENT 1���� (!AF_INE�pp�{�?!tcp{����!ud��ˎ!icm�����rkXY�Ӵ����q�)� p�/�A��p�)�j�M�Y���}��� �����ן���8�J� 1�n�U�����*�s����}}�����,�?,+��jfp�/z�֯�K�,������A��,  �p���@����ʿ�u"�ut�}��sF�P�PORT_WNUM�s�p��P�_CARTR�EP�p��|�SKS�TA�w K�LGmSm���������pUnothingϿ������c{t�TEMP �����ke��_a_seiban0C�, S�y�dߝ߈��߬��� ��	����?�*�c�N� ��r��������� ��)��M�8�q�\�n� �������������� #I4mX�|� �����3�ɟVERSI�p ��d disa�bled>SAV�E ��	2600H721:	&�!;���̏�� 	(�rmoN+E/`�eb/�/�/�/�/"�*z,�? %`����_-� 1���E0�b8eO?a?4g�npURGE_ENaB3��v�u�WF�0#DO�v��vWi��4��q*�WRUP_DELAY �C���5R_HOT �%�f�q:�.O�5R_?NORMALH
�xOrOAGSEMIQO�wO�OlqQSKIP-3���>3x$�O  _1_C_]&ot_b_�_ �_�_�_�_�_�_o(o :o o^oLo�o�o�olo �o�o�o $�oH 6X~��h�� �����D�2�h��z�����$RBT�IF�4G�RCVT�MOU\������DCR-3��I� �QE=U�4�1D͛�C��JA?͜6��ט]���q��6��1B��AY�����_V�R_ ;�x�5;��0;�i�;�du;�t�<!��h��R���̝�����&� 8�J�\�n�����������RDIO_TYPE  4=��¯�EFPOS1 1�C�
 x/:�H2 ��b�M���/��E�ο i�˿ϟ�(�ÿL�� pς��/�i��ϵ��� ��߭�6���3�l�� ��+ߴ�O����߅ߗ� ��2��V���z��� 9����o������� @�R�����9�������~�OS2 1��;+�u���-��Q���3 1������G���gS4 1�~���ZE|~�S5 1��%7q��/�S6 1Ũ��/��/o/�/&/S7 1�=/O/a/�/??=?>�/S8 1��/�/��/0?�?�?�?P?SM�ASK 1�߯ p)�OF�7XNOܯ�FUO_C�MOT�E���X4uA_CFG �|M�1\A�PL_RANGxA����AOWER ����@�FSM_�DRYPRG �%�%y?!_�ETA�RT ��N/ZU?ME_PRO�O_��_X4_EXEC_?ENB  ����GSPDdP�P�X��νVTDB�_�ZRM��_�XIA_OPT'IONφ����pAINGVERS.a��z_�)I_AIRPUR�@� @O�o�=MT_��0T�@zO��OB�OT_ISOLC�=N�F�1�a�eN�AMERl�bo�:O�B_ORD_NU�M ?�H�a�H721  �V1wLqr�qqrV0qr��s�ps�u\@��PC_OTIMĖ��x��oS232�B1�����aLTEAC�H PENDAN΀�7\H��x?c��Mainten�ance Con%sV2�#�"�_�No Use�� N��r���������С��rNPO>P�r\Az<e�qCH_LgP3�|Nw�	<��?!UD1:b�	�=R�0VAILRq2e���upASR  ��:a�B�R_INTVAL1f���I�+n��V_�DATA_GRP� 2���qs0DҐP�?`��?��o�� ������կï���� �-�/�A�w�e����� �����ѿ���=� +�a�Oυ�sϕϗϩ� �������'��K�9� [߁�oߥߓ��߷��� �������G�5�k�Y� ��}���������� ��1��U�C�e�g�y� ������������	�+Q?uDA�$S�AF_DO_PULS�pE@�C�� 'CAN�r1f�vp�SC�@�'��'Ƙ�Q+V0D�D�q(L�L�+AV2 y�' 9K]o���`����ڈ�%�2($Md($C!qu�1#
) @�C@o/�/�/�.W)k/ M���$�_ @݃T:`�/??&?39?T D��3?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|Ox֏��i%�O��O�O܉�!L� �;��o݄�p�M
�t��Dipp��L��J� � ��jL���j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����������(�:��� �/c�u���������Ϗ ��B�%�1�C�U� g�y���������Ƒ��0RMS�EW]�$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ�����M� ��*�<�N�`�r߄� �ߨ���������� &�8�J�\�ǟ����� ������������� ,�>�P�b�p������� ��������%7 I[m���� ���!3EWit�OB3t� ����////A/ S/e/w/�/�/�/�/�/��*��/?6���\R?�M	12345678XR�h!B!�)�����? �?�?�?�?�?�?OO A�>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_o]-O�_�_�_ �_�_�_�_o"o4oFo�Xojo|o�o�o�oq_BH�o�o�o!3 EWi{���������v[;�j�A�S�e�w����� ����я�����+�0=�O�a�xYD�k��� ����ɟ۟����#� 5�G�Y�k�}������� v_ׯ�����1�C� U�g�y���������ӿ ���	�ȯ-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�σ� �ߧ߹��������� %�7�I�[�m����D��v6����z���!�3�O:Cz � A�z   Ո@�2�v0� �@�
���  	�r�������������ph�u��� ��K]o���� ����#5G Yk}��0�� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-?G�������*@�  <X4t��$S�CR_GRP 1��'� '��� �t �t�� E5	 _�1��2 �2�4��W1G3�;97�7p�?�?OC��|�~BD�` D��3NGK)R-�2000iC/1�65F 5678�90��E��R�C65 �@�
O1234�E�6t�"A�����C�1F@�1�3�1)�1A�:�1�I	��?_Q_c_u_��_���H��0 T�7�2�_�?�_ �_o�6�t��_Lo��_poB8boK�h�@��UO��  uP��1BǙ�B�  B�33Bƿ`��e�b�c�1Ag��o # @t��e�1@>@	O  ?�w�bH�`�2�j�1F@ F�`\rd[o�s� ������*��9 �a�a)rU�@�R�d�v�B����ʏ���ُ ����H�3�l�W��� {���Ě2C�?����7���9�t�!q@"p>SԪD_�U�rh�`y��`ȏ��G �L�3��ϯ�A>G�1H��"oe��)�t� �<�N�\�*�pq�}���^� P���(����ӿ�g1EL�_DEFAULT�  �D���t���HOT�STR� ��MI�POWERFL � K����?�WF�DO� S�RV�ENT 1�����P0� L!DUM_EIP�����j!AF_�INE��ϵ!�FT�������!��_B� ��i�!�RPC_MAI�Nj�LغXߵ�|�V�IS��Kٻ���!7TP��PU�߳��d��M�!
PMON_PROXYN�e<���g��f�����!RDM_'SRV���g��1�G!R�DM���h ��}�!
~�M���i�l���!RLSY1N�@����8���!ROS��<�y4a!
CE��MTCOMb��k�P�!	vCON�S���l��!>vWASRC ����m�E!vUS	BF��n4�0ߵ ����/�'/��K//o/�RVICE_KL ?%��� (%SVC�PRG1v/�*�%2��/�/� 3�/�/� 4�??� 56?;?� 6^?c?� 7�?�?� \�$�?L19�?�;�$H� O�!�/+O�!�/SO�!  ?{O�!(?�O�!P?�O �!x?�O�!�?_�!�? C_�!�?k_�!O�_�! AO�_�!iO�_�!�Oo �!�O3o�!�O[o�!	_ �o�!1_�o�!Y_�o�! �_�o�!�_{/�"� �/ � F�E1���� ����
�C�U�@� y�d����������Џ ����?�*�c�N��� r��������̟�� )��M�8�_���n��� ��˯���گ�%�� I�4�m�X���|������ǿ�ֿρ*_DE�V ����MC:�H'�GRP 2ׇ�+p� �bx 	� 
 ,y�ϒ�+r ~ϻϢ���������� 9� �]�o�Vߓ�z߷� �߰������#�z�G� ��k�}�d������� ���������U�<� y�`���������*��� 	��-QcJ� n����� �;"_FX��� �����/�/ I/0/m/T/�/�/�/�/ �/�/�/�/!??E?W? �{?2?�?�?�?�?�? �?O�?/OOSO:OLO �OpO�O�O�O�O�O_ ^?�O=_�Oa_H_�_�_ ~_�_�_�_�_�_o�_ 9oKo2oooVo�ozo�o �o _�o�o�o#
G .@}d���� ����1��U�<� y����o��f�ӏ�̏ 	���-�?�&�c�J��� n��������ȟ�� ��;���0�q�(���|� ��˯���֯�%�� I�0�m��f�����ǿp������R�d ��	�4��X�C�|�gό�ϯ�%�����R������������� ��+��O�=�s߁��� ����i���������� 	��Q��x��A�� ����������Y�� P���)���q������� ����1�U���I�� Ym���	� -�!E3U{ i������ //A///Q/w/��/ �g/�/�/�/�/?? =?/d?v?-?O?)?�? �?�?�?�?OW?<O{? OoO]OO�O�O�O�O �O/O_SO�OG_5_k_ Y_{_}_�_�__�_+_ �_ooCo1ogoUowo �_�_�oo�o�o�o 	?-c�o��oS �O�����;� }b��+��������� ɏ�ݏ�U�:�y�� m�[��������ş� -��Q�۟E�3�i�W� ��{����دꯡ�ï ���A�/�e�S���˯ ���y��ѿ���� =�+�aϣ���ǿQϻ� �����������9�{� `ߟ�)ߓ߁߷ߥ��� ����A�g�8�w��k� Y��}�������� =���1���A�g�U��� y����������	�� -=cQ���� ��w���) 9_���O�� ��/�%/gL/^/ /7///�/�/�/�/ �/?/$?c/�/W?E?g? i?{?�?�?�??�?;? �?/OOSOAOcOeOwO �O�?�OO�O_�O+_ _O_=___�O�O�_�O �_�_�_o�_'ooKo �_ro�_;o�o7o�o�o �o�o�o#eoJ�o }k������ ="�a�U�C�y�g� ������ӏ���9�Ï -��Q�?�u�c���ۏ ��ҟ�������)�� M�;�q�����ןa�˯ ��ۯݯ�%��I��� p���9�����ǿ��׿ ٿ�!�c�Hχ��{� iϟύ��ϱ���)�O�  �_���S�A�w�eߛ� �߿����%߯��� )�O�=�s�a���߾� �߇�������%�K� 9�o������_����� ������!G��n ��7������ O4F��g �����'/K �?/-/O/Q/c/�/�/ �/��/#/�/??;? )?K?M?_?�?�/�?�/ �?�?�?OO7O%OGO �?�?�O�?mO�O�O�O �O_�O3_uOZ_�O#_ �__�_�_�_�_�_o M_2oq_�_eoSo�owo �o�o�o�o%o
Io�o =+aO�s�� �o�!���9�'� ]�K��������q��� m�ۏ���5�#�Y��� ����I�����ßşן ���1�s�X���!��� y���������ӯ	�K� 0�o���c�Q���u��� �����7��G��;� )�_�Mσ�qϧ���� ϗ�ߓ��7�%�[� I���Ϧ���o����� �����3�!�W��~� ��G����������� 	�/�q�V������w� ����������7�. ����O�s�� ��3�'7 9K�o��� ���#//3/5/G/ }/��/�m/�/�/�/ �/??/?�/�/|?�/ U?�?�?�?�?�?�?O ]?BO�?OuOO�O�O �O�O�O�O5O_YO�O M_;_q___�_�_�_�_ _�_1_�_%ooIo7o mo[o}o�o�_�o	o�o �o�o!E3i�o ��Y{U��� ��A��h��1��� ������������[� @��	�s�a������� �����3��W��K� 9�o�]���������� �/�ɯ#��G�5�k� Y���ѯ������{� ����C�1�gϩ��� ͿW��ϯ�������� 	�?߁�fߥ�/ߙ߇� �߫��������Y�>� }��q�_����� �����������7� m�[����������� ����!3iW ������}�� �/e��� U����/�/ m�d/�=/�/�/�/ �/�/�/?E/*?i/�/ ]?�/m?�?�?�?�?�? ?OA?�?5O#OYOGO iO�O}O�O�?�OO�O _�O1__U_C_e_�_ �O�_�O{_�_�_	o�_ -ooQo�_xo�oAoco =o�o�o�o�o)ko P�o�q��� ���C(�g�[� I��m�������ُ�  �?�ɏ3�!�W�E�{� i�����؟���� ��/��S�A�w����� ݟg�ѯc�����+� �O���v���?����� Ϳ��ݿ��'�i�N� ��ρ�oϥϓ��Ϸ� ����A�&�e���Y�G� }�kߡߏ�������� ���߱��U�C�y�g�����������$S�ERV_MAILW  �����OUTPUT����RV 2�v��  � (��x��_���SAVE����TOP10 2}�9� d 	� ��������+= Oas����� ��'9K] o������� �/#/5/G/Y/k/}/`�/�/�/���YP|����FZN_CFGw ڍ����j��!GRP �2��'&� ,B�   A=0��D;� B>0�  �B4��RB2�1l�HELL�"!܍�$�L�M�7�?>�;%RSR�?�? �?O�?%OOIO4OmO XOjO�O�O�O�O�O�O�_!_3^�  ��R3_a_s_AR_ ���{_�R�P�xWIR2��d�\�]�R�h6HK 1�v; �_o"ooFooo jo|o�o�o�o�o�o�o �oGBTfb<?OMM �v?��g2FTOV_EN�B��A�$��ROW_?REG_UI����IMIOFWDL�pߥ~@5�WAIT�r�Y�8���v�@�0�TIM�u��j�VA��A��_UNIT�s��$��LC�pTRY�w�$���MON_ALIAS ?e�yH�he��%�7�I� [�i��������m� ���
��.�ٟR�d� v�����E���Я��� ���*�<�N�`��q� ������̿w���� &�8��\�nπϒϤ� O���������߻�4� F�X�j�ߎߠ߲��� �߁�����0�B��� f�x����Y����� ������>�P�b�t� ������������� (:L��p�� ��c�� � 6HZl~)�� ����/ /2/D/ V//z/�/�/�/[/�/ �/�/
??�/@?R?d? v?�?3?�?�?�?�?�? �?O*O<ONO`OO�O �O�O�OeO�O�O__ &_�OJ_\_n_�_�_=_ �_�_�_�_�_�_"o4o FoXooio�o�o�o�o oo�o�o0�oT fx��G��� ���,�>�P�b�� ��������Ώy�����(�:���$SM�ON_DEFPR�O ����c� �*SYSTEM*�M�RECALL �?}c� ( ��}4xcopy �fra:\*.*� virt:\t�mpback��=�>192.168�.56.1:11620 ԑ۟�����}8��s:or�derfil.dat��ßٟj�|���{}/��mdb:���G�ՐS������3 ������Еׯh�z��� ���3�E�X������ }
xyzra?te 61 ���� ҿc�uχ��#�C�7188 A�S��������tpdiosc 0��8 �����b�t߆��tpconn 0 ,�@>�P�������7#��5�+�8�k�}��. ��>��R�������2#�6ϲ���g�y��� ���<���W����� �1����fx��� 8��S���� ��Q�bt�����<�����/�e 1�,Ͼ�a/s/�/�0��:pickupw.tp1%emp����U/�/�/
?��:place�/J�/e?w?�?��@? �?S?�? �?O/�߿?�?bOtO �O�?�?=OOO�O�O_ O)O�O�O^_p_�_�O �O9_K_�_�_ o_%_ �_�_Zolo~o�_�_5o GoYo�o�o!o�o�o �ohz��o1CU`��
���{36U� ��e�w����0�?� Q������-}��͏ ^�p����/�/8?8�T� ���	�?.?��R�c� u���,�H�ۯ� ������7�үc�u� ���?/;�V���� Ϟ����ѐ׿h�z� �ϟ���:�U�����
� ���A���d�v߈ߚ���$SNPX_A�SG 2�������� �>���%����� � ?���PARAoM ���ѯ �	��P�������*����O�FT_KB_CF�G  �ô՞�O�PIN_SIM + ��%��������RVQST_P_DSBk�%�|���SR ��� � & C�ONROD��/����TOP_ON_ERR  /��W�L�PTN z���AH��RING_PRM�V� ��VCNT?_GP 2��'���x 	��������� ��$��VD��ROP 1���(� ��_q���� ���%7I [m������ ��/!/3/Z/W/i/ {/�/�/�/�/�/�/�/  ??/?A?S?e?w?�? �?�?�?�?�?�?OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_r_o_�_�_�_�_�_ �_�_�_o8o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy �������	� �-�?�Q�c������� ����Ϗ����)� P�M�_�q��������� ˟ݟ���%�7�I� [�m��������ܯٯ�����!�3�=PRG_COUNTL����[�_�ENBĔ�Z�M��N䑿_U�PD 1��T  
H���ۿ��� (�#�5�G�p�k�}Ϗ� �ϳ����� ����� H�C�U�gߐߋߝ߯� �������� ��-�?� h�c�u������� ������@�;�M�_� ���������������� %7`[m ������� 83EW�{�� ����///// X/S/e/w/�/�/�/�/ �/�/�/?0?+?=?O?�x?s?�?Q�_INF�O 1�ɹ�� ��F��?�?�?O�9��]MEA?�>�>�O�7���PA6�SB���u�P�YS�DEBUGi�ʰ��0d��z@SP_PwASSi�B?�K�LOG �ɵ����0>H�? � ����1UD�1:\�D�>�B_M�PC�Mɵ:_L_ɱ��Aj_ ɱVSAV ��MA�A�B�5� XSVnKTE�M_TIME 1u��G�� 0�0��4�lXl_�0���T1SVGUNS�İj�'���`A�SK_OPTIO�Ni�ɵ����?a_�DI�@��[eBC2_GRP 2�ɹ��U�o�0@�  C���cP��`CFG 3�k�\ �V�f`
EOB-R xc������ ���>�)�b�M��� q���������ˏ�� (��L�7�p����Vn� ��n�ϟ�\����� ;�&�_�q^�QdT��� ����ѯ������� )�+�=�s�a������� ��߿Ϳ���9�'� ]�Kρ�oϑϓϥ��� �Ȭ�����1�C��� g�U�wߝߋ������� ��	���-��Q�?�a� c�u���������� ��'�M�;�q�_��� ������������ 7��Oa��! �����!3E iW�{��� ��/�///S/A/ w/e/�/�/�/�/�/�/ �/??)?+?=?s?a? �?M�?�?�?�?O�? 'OO7O]OKO�O�O�O sO�O�O�O�O_�O!_ #_5_k_Y_�_}_�_�_ �_�_�_o�_1ooUo Coyogo�o�o�o�o�o �o�?!?Qc�o �u������ �)��M�;�q�_��� ����ˏ���ݏ�� 7�%�G�m�[������ ��ٟǟ����3�!� W�o�������ïA� �կ����A�S�e� 3���w�����ѿ��� ���+��O�=�s�a� �υϧ��ϻ������ �9�'�I�K�]ߓ߁� ��m��������#�� G�5�W�}�k����� ���������1��A� C�U���y��������� ����-Q?u c������� ��/A_q� �����/� ��$TBCSG_�GRP 2����  ��  
 ?�  J/\/F/�/j/�/ �/�/�/�/�/;#"*#��1,d0�?1?!	 HD� 6s33[23�\5O1B�!x?ޅ9D)�6L�=ͣ1>���g6�0�CF�?�?�8fff��1�>��!OICj˱�6�1H4B��C{OO)H�d�0|A�]0@HDO _O)H�1�8CFr�O�M@ �. XU&_�O_�Q_n_9_K_�_�_�[?��0�Sp �	�V3.00�R	�rc65�S	* `�T"o�V|A�0 58 `�Y G`m�Ho  � �%@��_�o�c#!J2*#��1-�o�hCFG ��;!C!�j��B"]b�l|�BPz�Pv a������� ��<�'�`�K���o� ������ޏɏ��&� �J�5�n�Y�k����� ȟ������\	�� -�ן`�K�p������� ��ޯɯ��&�8�� \�G���k�����!/ ۿ�����5�#�Y� G�}�kϡϏϱ����� ������C�1�S�U� gߝߋ��߯�����	� ���?�-�c�Q��� Y����m������)� �M�;�q�_������� ����������%I [m9���� ���!E3i W�{����� /�///?/A/S/�/ w/�/�/�/�/�/�/? +?��C?U?g??�?�? �?�?�?�?�?OO9O KO]OoO-O�O�O�O�O �O�O�O_�O!_G_5_ k_Y_�_}_�_�_�_�_ �_o�_1ooUoCoyo go�o�o�o�o�o�o�o 	+-?uc� ���y?���� ;�)�_�M���q����� ��ݏ�����7�%� [�I��������o�ٟ ǟ����3�!�W�E� {�i���������ï�� ���A�/�e�S�u� ���������ѿ��� ��+�a��yϋϝ� G��ϻ������'�� K�9�o߁ߓߥ�c��� ��������#�5�G�� �}�k�������� ������C�1�g�U� ��y�����������	 ��-Q?a�u ������� /���q_��� ����/%/7/� /m/[/�//�/�/�/ �/�/?�/?!?3?i? W?�?{?�?�?�?�?�? O�?/OOSOAOwOeO �O�O�O�O�O�O�O_ _=_+_M_s_a_�_ C�_�_}_�_�_o9o 'o]oKo�ooo�o�o�o �o�o�o�o#Y k}�I���� �����U�C�y� g���������я��� �	�?�-�c�Q�s�u� �������ϟ��)� ;��_S�e�w�!����� ˯��ۯݯ�%��I� [�m��=�����ǿ����վ  ��� �)���$T�BJOP_GRP� 2�ݵ�  ?��i	A�H��O���� ��ߐpXd� ����� � �{,� @��`�	 �D ���CaD�q��`���fff���>��H�ϻ�L̽�	�<!a���>����=�B� � Bp��8�C�D�)�U�CQp�Dw�S�Ι��yҜ��v� ?�����?�\<���U�ҷ��%�CV+��x/���S�D5mi��{Բ��ع�<����z�>\>��33C�  CqA��`�K�j��u��bߐ���z�;�9�bB�E�>���׵ҳ� C��V���s����&��ǌ?��;��6��%�~]�D&� C����������
Ѷ� ?�s33����<Z;]u���ff�ҴK������U�)C- _i�u���� ��*IcM������Ƙ�����	V3.00�f�rc65e��* e��/ ' �F�  F��� F� F� � G� GX� G'� G;�� GR� Gj`� G�� G�|� G� G��� G�8 G��� G�< H� H� H���2 Ez  E�@� E�� EB F� FR FZ F��� F� F�P�<"G � Gp�L#?h GV� �GnH G�� �G�� G�( �=u=+*�(�$`Q�?�2�3?� � ��M?[:A��*�SYSTEM
!V�8.30218 ��38/1/201�7 A y  �p7M�TP_T�HR_TABLE�   $ $�1ENB��$D�I_NO��$D�O�4  ��1C�FG_T  �0�0MAX_IO�_SCAN�2MI�N�2_TI�2DM�E\��0@�0 � � $CO�MMENT �$CVAL	CT~�0PT_IDX��uEBL�0NUMQB�ENDIJfAZITI�D]B $DU�MMY13��$�PS_OVERF�LOW�$�F��0FLA�0YPE��2�BNC$GLB_TM�7�EF@�1�0ORQCTRL�1��$DEBU�G�CRP�@2@ � $SBR_P�AM21_VP� T$SV_ER�R_MODU4SC�L�@RACTIO��2�0GL_VIE�W�0 4 ]$PA$YtRZtR�WSPtR�A$C�A@A�6aQUeU� �0N�P3@$�GIF3@}$eQ �lP_S�PiQ L�pP�VI<P�PF�RE��VNEARPLA�N�A$F	iDI�STANCb�1J�OG_RADiQ�@$JOINT�SP尤TMSE]TiQ  �WE�UACONS2@B�R�ONFiQ	� �$MOU1A`��$LOCK_FOyL�A�2BGLV@C�GL�hTEST_sXM@@raEMPE`�,R�b�B`�$U1S;AfPH`2P�S:�a�bMP_�`�a=QCENEdRr� $KARE�@M>�3TPDRAhP;t>2aVECLE�32dkIU�aqHE�`�TOOLH`�0qsV�I{sRESpIS3�2�y64�3ACH4X`�`~qONLE�D�29�B�pI�1 � @$RAIL__BOXEHaPoROBO�d?�Q?HOWWAR�0�r<�@�qROLM�B�A�C �SK�r�@�07O_F9�!��St�qiQ
>o �RVp�OCiQ_�SLO�GaK��VOUZb�R�eAELEC�TE<P`�$PI=P�fNODE�r�r��qIN�q2^��pCORDED�`�`}��0P9P@  wD �@OBAU`TA�a����C�@��p�P�q0��ADRAܥ0F@TCHup 7 ,�0EN�2�1A�a_�Tl�Z@�BޣRVWVA!A� � ApeR�5P�REV_RT�1�$EDIT��VS�HWR9�S@	UАI�S`yQ$IND�0@1QB蓗q$HEAD�5@ ��p5@溒KEyQ�@CPS�PD�JMP�L��5�0RACE�4U�a�It0S�?CHANNEzp��	WTICK{s�1M�`A�0@�HN�A�D0^�]D�`CG�P8���v�0STYf��q�LO�A�3B���jP� t 
��Gr�%�$���T=PS�!$UNIGa5A�E��0�FPORT��SCQU5ptR���B��TERCJ@���T=SG� �PPL6�$�DE��$`Thqb�0OK@>CV�IZ�D4�Q�E�APR�A�Ͳ�1��PU}aݵ_�DObk�XSV`KN�6AXI��7�qgUR_s�E$T�p���*��0FREQ_,hp<�ET=�P�b�OPARA`@.P
@�:[���ATHr�3@a�D�s�s�0 �2�SR_Q�0l8}��@�1TRQIc���$`�@��BRup��VyE@@��NOLD��AAp7a��x@�A��AV_MG����¨/���/�D)�D;�D�M�J_ACC.�C��<�CM��0CYC0M@3@��M@_E������٘@NbSSC��@  hPD1S���1�@SP�0*�AT:����@��i��B�ADDRES{sB���SHIF}b�a_W2CH�@&�I�@�|��TV�bI�2�]��h>��C�
�j
��2V����0 \��������웱�@��CnӞ�aºꯆ:R����TXSCREE���0�TIN!AWS�P;��T0r�sQ_>�jP TQ� 7P�B�6QP��
���
���RROR_�"a�@���E�UE�G� ���U��@S�XQ�RSM�� �U�NEXg��6��0S_�S��	0���>�C�b��o� 2m6�UE���2�GRUͰGMTN_KFLQ�#POHg/BBL_�pWg@�0� ����O�QƾLEn���pTO�`C�RIGH�B�RDITd�CKGRg@�TEX,���WIDTH�sݐBh�A�A{q��I_/@�H��  8 $LT_ �|�Y0@RyP�b�s�w�B��RGOu��0D0TW�� U� �R�b�L�UM�!�^�ERV���]PFP`>��1z'@r�GEUR�ciF\��Q)��LP�Z�Ed��)'�$(P�$(�p#)5!+6!+7!+8"b�>CȰ`���F�q�aS�@�EUSReT  <��/@U�R��R�FOChq�PPRI�z�m�@?A� TRI}P�qm�UN�0
�4!�P ��0�5�p7��b;�5� "T\� ̱G �T7����}�O2OSNAd6R A���;3wq�1#n_�S �^�2�����aU!"A�$�?�?+"��;3OSFF�` P%O��3=O@ 1#PD:,D$PGUN#K`}S�B_SUBB�Pk SRT�0��&0��"avp��OR�p�E'RAU���DT�Ib���VCC��H�' ���C36MFB�1ĢSPG?�(s (b`�STE�Qaʀ9PWTѠPE�:��GXd) ����J�MOVE��{Q6RA�N4`?[�3DV�S6RLIM_X�3qV�3qV \XvQk\:V1�IP&�2VF��C砽@d��G�*��IB�P,�S� _�`�p�b����@ (0G�B�� "P�@��pr+�x �r �,� tRn@��s C@TeGDRI�PSfQV!��wdԐ��D�$MY_UBY�$\d�;QA��S���h�q�bP_�S�ף�bL�BMvkQ$j�DEYg��EX� ���BUM_�MU6�X�D<q U�S�?��;VGo�PACI�TP�<Uyr��3yrkSyr:;qRE0nr�1l�9cyrz�@,�BTARGP!P�p�R<aR{0�@�- d��;cB	4:r��R�DSWqp�S�n�:s˰O�!d�A(v�3���E��U�p0Zm��vHK�.���K�AQ��0���?SE9A����WOR�@3���uMRCVr/ U��O��M�@C��	ÂC�sÂREF ��̆��gRj�
��  Ȋ�ي��=�̆r�_RC��s�����@`����b������to0 �Т�;��4� �e�OU���rH��\c(`+�u��2��0<���̰� -=��Ѻf�K�SUL3a.2�C7Po/+p�NT�a��]��ag��g��!g�&�L�c���cP������!�@T���s�1���o@APg_HUR�ۥSA>SCMP��F����
�_&�R�T�����X.���VGFS��E2d �M8� � Y0UF_�����J��RO� ���l�W,rUR�GR�mq�I���D_V_h[�D�@zY��3�WIN".rH���X-V
A�RqR�P�WEw�w�q`|c6v,q��RvLOiP�tc�PMc��3t� +=�PA' =�CACH6�����@��,p����K�ۓC�Q-Io�FR"�T� $�N��$HO�@�R�� `�rc��[�֘p���ڔ�VP�r����_'SZ3p���6����12� ��]p�؆P�؛WA3�MP��aIkMGx���AD鞨qIMREٔ6�_SIZ�P��!po��6vASYNBUF6vVRTDh�t�F�~OLE_2D�T(��t��0C0aUs��yQP�X�ECCU�x�VEM�p����#�V�IRC��VTP �����G�p��t��LA�s�!���Mco�4��;�CKLA�SQC	��ђ�@5 ! �A�� @&B�Tq$��$`��6 |F@o���Xñ�T�o�?a��"�uI���r/��`�BG� VEJ�`P�K|p1���֖K�MH�O+��R7 � �}F���ESLO�W}w]RO>SAC�CE*@-�=�xVR`:��11�yrAD��/0rPA��&�D:�1�M_Ba�81N��JMP���A8y�>b�$SSC6u���M��C��@92��S�8��N/�PLEX���: T〲C�Q���6�FLD?1DEZ�FIQ rO�qt�y� K�P2��;O� ϱPV�>��MV_PIZ���G�BP��`а�FIQ�PZ�$���0����GA%p��LOO0Tp�JCB�T*����� ��ړPLCAN�R&�L�F�� �cDV�'M�p���U�$�S�P.q�%�!��%#�㱶C4G�����RKE�1�V�ANC]K�A0p K<�@�?�?Q3A�a =�?q??Tp0�9����r> hܰ��	��K9�fA2b<LX@̠OUe�ݒA��Y
O���SK(�M��VIE�p2= pS0:�|R? <{@xX���`UMMY�����Re��D��MȧCU�`b�U�@�@ $�@TIT> 1$PR8�U�OPT�VSH�IFʀ�A`��a���D�0����$�_R$�UړQ.q Z�U�s�ot�QavȆQ5fSTG@cVSC9O��vQCNT���3 � }w�RlW�RzV�R�W@�R�XLo^opjjA2���51D>a�0� ]�pSMO��B%dTC�J�@1u���I_���@C%�Gi��LI� '��XV�R�DDY�@T���ZABCP��E�r�b���
J�Z�IP�EF%��LVҡ�L����ZM�PCF�eGy�$�p	�rDMY_�LN$@Ar8��dH� ���g��>�MC�MİC��CART�_Xq�P�1 '$JvsptD��|r��r�w���u���UX�W�puUXEUL�x�q�u�t�u�q�q��y�q�v r�eI �Hk�d���Y�`D>�� J 8o�	V��EIGH��H?�("��f��ĔK� �= �C���`$B&�K���1_�B��Lg�RV� F�`��COVC؀qrfq9��@}�De�
����7�D��TRȰ	�V�1�S3PH� ǑL !�S��i�{����ST�S  ��������u�<�ѐNa�1 ����C �������������������U����	��
��Q����������p����( ��RDI������ğ֟����t�O|���������ί$ஔ�Sz��� >��� ��ſ׿�����1� C�U�g�yϋϝϯ��� �������v�}���8� !�3�E�W���'�9�`K�]���� �����U��� p��( ��� ���@A�v�^`BF_�TT��ի���I�V�>0n�J�_�I�R {1&� 8��Ȩ�%к� ��C�   ������������"� 4�F�X�j�|������� ������1gB Tjx���� �р����0B QI�ZlJ� ��������/ "/4/F/X/FҒ�t/�/�b*���/�/��bv�@�`�v�MI_CH+ANU� `� #3�dbV�`�u�&0ET>�_AD ?��y0�m��/�/�?�?زd0RLPs�!&�!��4�?�<SNMA�SKn8��1255.4E0�33OEOWO~�OOLOFS^Q�  �%X9ORQCTRL &�"V�m��O��T�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo�(l�OKo:ooo��PEΌpTAIL8�JPG�L_CONFIG� 	�ᄀ�/cell/$C�ID$/grp1�so�o�o1�#� �?\n����E ����"�4��X� j�|�������A�S�� ����0�B�яf�x� ��������O����� �,�>�͟ߟt���������ίB�}c��� (�:�L�^���`o��e��b���Ϳ߿��� \�9�K�]�oρϓ�"� �����������#߲� G�Y�k�}ߏߡ�0��� ���������C�U� g�y����>����� ��	��-���Q�c�u� ������:������� );��_q�� ��H��% 7�[m�����]`�User View �i�}}1234567890�
//./�@/R/Z$� �cz/���2�W�/�/�/�/ ??u/�/�3�/d? v?�?�?�?�??�?�.4S?O*O<ONO`OrO�?�O�.5O�O�O�O@__&_�OG_�.6�O �_�_�_�_�_�_9_�_�.7o_4oFoXojo|o�o�_�o�.8#o�o�o�0B�ocir �lCamera��o������NE�,�>� P��j�|�������ď�I  �v�)��&� 8�J�\�n�������� �ڟ����"�4�[��vR9˟�������� ȯگ�����"�m�F� X�j�|�����G�Y�I 7�����"�4�F�� j�|ώ�ٿ�������� ��߳�Y�����Z�l� ~ߐߢߴ�[������� G� �2�D�V�h�z�!� �unY���������� ���B�T�f������ ����������Y�"i{� 0BTfx�1�� ���,> P��Y��i���� ����/,/>/� b/t/�/�/�/�/cu9H/�/?!?3?E?W? �h?�?�?F/�?�?�?��?OO/O�j	�u0 �?jO|O�O�O�O�Ok? �O�O_�?0_B_T_f_ x_�_1OCO�p�{._�_ �_oo+o=o�Oaoso �o�_�o�o�o�o�o �_�u���oOas� ��Po���<� '�9�K�]�o�PEc� ���͏ߏ���� 9�K�]����������� ɟ۟����ϻr�'�9� K�]�o���(�����ɯ �����#�5�G�� ��;�ޯ������ɿۿ ���#�5π�Y�k� }Ϗϡϳ�Z�����J� ���#�5�G�Y� �}� �ߡ������������<���  ��N� `�r���������x����   $� ,�J�\�n��������� ��������"4F Xj|����� ��0BTf x������� //,/>/P/b/t/�/��  
��(  ��B�( 	  �/�/�/�/�/??8? &?H?J?\?�?�?�?�?t�?�*4� �n� O1OCO��gOyO�O�O �O�O��O�O�O_VO 3_E_W_i_{_�_�O�_ �_�__�_oo/oAo So�_wo�o�o�_�o�o �o�o`oroOa s�o������ 8�'�9��]�o��� �������ۏ���F� #�5�G�Y�k�}�ď֏ ��şן�����1� C�U���y�������� ӯ���	��b�?�Q� c�����������Ͽ� (�:��)�;ς�_�q� �ϕϧϹ� ������ H�%�7�I�[�m���� �ߵ���������!� 3�E�ߞ�{����� ����������d�A� S�e������������ ��*�+r�Oa�s������0@ A�������� ��)frh:�\tpgl\ro�bots\r20�00ic6_16?5f.xml�` r�������/����/3/E/W/ i/{/�/�/�/�/�/�/ �//
?/?A?S?e?w? �?�?�?�?�?�?�?? O+O=OOOaOsO�O�O �O�O�O�O�OO_'_ 9_K_]_o_�_�_�_�_ �_�_�__�_#o5oGo Yoko}o�o�o�o�o�o �o o�o1CUg y�������o ��-�?�Q�c�u����������Ϗ���K � 88�?��2�� .�P�R�d��������� �П���(�R�<��^���r�����ܫ�$�TPGL_OUT?PUT ����_ ��� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ������ˠ2345?678901���� ����0�8�����_� q߃ߕߧ߹�Q߽��� ��%�7���}A�i� {����I�[����� ��/�A���O�w��� ������W����� +=����s��� ��e�'9 K�Y����� as�/#/5/G/Y/ �g/�/�/�/�/�/o/ �/??1?C?U?�/�/ �?�?�?�?�?�?}?�? O-O?OQOcO�?qO�O@�O�O�O�OyO֡}��_)_;_M___q_�]@���_�_� ( 	 ���_�_o�_ 5o#oYoGoioko}o�o �o�o�o�o�o/ UCyg���������	�?��Ƭ �-�G�u���c����� ��ߏ���`��,�Ώ P�b�@��������Ο p�ޟ����:�L��� p���$�������ܯ� X���$�Ư�Z�l�J� �����ƿؿz���� �2�DϮ�0�zό�.� ���Ϡ�����b��.� ��R�d�B�tߚ��� ���߄�����<�N� ��r��&������ ��Z�l�&�8���\�n� L����������|��� �� FX��|� 0�����d 0� fxV�� ���//�>/ P/�</�/�/:/�/�/�/�/?
2�$TP�OFF_LIM �[��@W����A2N_SV#0 � �T5:P_M�ON S��74�@�@2�U1S�TRTCHK �S�56_=2VT?COMPATJ8�1�96VWVAR �j=�8N4 R�? O�@}21�_DEFPROG� %�:%CO�NROD&O�?_D?ISPLAY*0�>�?BINST_MSwK  �L {J?INUSER�?�D�LCK�L�KQUI�CKMEN�O�DS7CREPS��2?tpsc�D�A�1P6Y52GP_KYST��:59RACE_COFG �Fr1�4u.0	D
?��X�HNL 2�93��Q�; $B�_�_o� o2oDoVohozj�UI�TEM 2�[� �%$1234?567890�o�e  =<�o�o�os�  !{!@ �oZC�o{�o�� �9K�o/�� ?�e������#� ��G���+���O��� ŏ׏Q�����͟ߟC� �g�y����]����� �������-���Q�� u�5�G���]�ϯ!��� �ſ)�տ���q�� ������3�ݿ�ϯ��� %���I�[�m���	ߣ� c�u��ρ������3� ��W��)��?���� ���ߧ�����c�S� e�w������k��� �����+�=�O���s� EW��c���� ��9�o� �n�����# �G�"/}=/�M/ s/�/��///1/�/ U/?'?9?�/]?�/�/ �/i?�??�?�?Q?�? u?�?PO�?kO�?�O�O@O�O)O;O_�TS�R��_UJ�  ��bUJ �Q`_UI
� m_�_z_�_8Z�UD1:\�\���QR_GRP 1��k� 	 @`@o!koAo/oeoSo�own��`�o�j��a�_�o�o�e?�  '9{#YG} k������� ��C�1�g�U�w����	�E��ÏSSC�B 2%[  �!�3�E�W�i�{������\V_CON?FIG %]�Q�]_�_���OUTP�UT %Y�����S�e�w��� ������ѯ����� +�_A@�S�e�w����� ����ѿ�����+� <�O�a�sυϗϩϻ� ��������'�8�K� ]�o߁ߓߥ߷����� �����#�5�F�Y�k� }������������ ��1�B�U�g�y��� ������������	 ->�Qcu��� ����); L_q����� ��//%/7/H[/ m//�/�/�/�/�/�/ �/?!?3?D/W?i?{? �?�?�?�?�?�?�?O O/OAOݟ�>�O�O �O�O�O�O�O�O_!_ 3_E_W_J?{_�_�_�_ �_�_�_�_oo/oAo Sod_wo�o�o�o�o�o �o�o+=Oa ro������� ��'�9�K�]�n�� ������ɏۏ���� #�5�G�Y�j�}����� ��şן�����1� C�U�g�x��������� ӯ���	��-�?�Q� c�t���������Ͽ� ���)�;�M�_�p� �ϕϧϹ�������� �%�7�I�[�m�~ϑ� �ߵ����������!��3�E�W�i�LH�������s���hO ������1�C�U�g� y���������t����� 	-?Qcu� ������� );M_q��� ����//%/7/ I/[/m//�/�/�/�/ ��/�/?!?3?E?W? i?{?�?�?�?�?�?�/ �?OO/OAOSOeOwO �O�O�O�O�O�?�O_ _+_=_O_a_s_�_�_ �_�_�_�O�_oo'o 9oKo]ooo�o�o�o�o �o�o�_�o#5G Yk}����� �o���1�C�U�g��y���������ӏ����$TX_SCRE�EN 1��w���}��@&�8�J�\�n���� �����ҟ����� ����P�b�t������� !�ίE����(�:� L�ïp�篔�����ʿ ܿ�e�w�$�6�H�Z� l�~������������ ��� ߗ�D߻�h�z� �ߞ߰���9�K���
� �.�@�R���v��ߚ��������k����$UALRM_M_SG ?��� ��zJ�\����� ��������������/�"SFw+�SEV3  �E��)�ECFG ���  �u@�  A�   ;B��t
 x�s �0BTfx�������GR�P 2� 0��v	 �/+�I�_BBL_NOT�E �
T��l�r��q�� +"DEFPR�O5�%9� (% k�/�p�/�/�/�/�/ ?�/%??6?[?F??�j?�?!,INUSE�R  o-/�?I�_MENHIST� 18��  �( | ��(/�SOFTPART�/GENLINK�?current�=menupage,153,1�?0`OrO�O�O�)'O9N?381,23�O�O��O	_�O+�O9Eed�itEBCONRODMOi_{_�__�?�_ �_�_�_oo�_AoSo eowo�o�o*o�o�o�o �o�o�oOas ���8���� �'��8V""A�_�q� ���������ݏ�� �%�7�Ə[�m���� ����D�V�����!� 3�E�ԟi�{������� ïR������/�A� Я�w���������ѿ `�����+�=�O�:� L��ϗϩϻ������ ��'�9�K�]��ρ� �ߥ߷�������|�� #�5�G�Y�k��ߏ�� ��������x���1� C�U�g�y�������� ��������-?Q cu`�rϫ��� �);M_q ������/ /�7/I/[/m//�/  /�/�/�/�/�/?�/ 3?E?W?i?{?�?�?.? �?�?�?�?OO�?AO SOeOwO�O�O���O �O�O__+_.OO_a_ s_�_�_�_8_J_�_�_ oo'o9o�_]ooo�o �o�o�oFo�o�o�o #5�o�ok}�� ��T����1� C��g�y�����������O��$UI_P�ANEDATA �1������  	��}/frh/c�gtp/whol�edev.stm�ӏ1�C�U�g�R�)Gpri���]�}���Ɵ؟���� � ) "�F�-�j�Q������� į��������B�pT�;�x�V���A������Ŀֿ��� �_�0ϣ�B�f�xϊ� �Ϯ���'�������� �>�%�b�I߆ߘ�߀�ߣ�������  ��8���T�Y�k�}�� ������J����� 1�C�U���y���r��� ��������	��- QcJ�n��0� B��);M� q������� /h%//I/0/m// f/�/�/�/�/�/�/�/ !?3??W?���?�? �?�?�?�?:?OO� AOSOeOwO�O�OO�O �O�O�O�O_ _=_O_ 6_s_Z_�_�_�_�_�_ �_d?v?4O9oKo]ooo �o�o�_�o*O�o�o�o #5�oYkR� v������� 1�C�*�g�N�����o "oӏ���	��-��� Q��ou���������ϟ �H���)��M�_� F���j�������ݯį ����7�����m�� ������ǿ����p� !�3�E�W�i�{�⿟� �����ϼ������/� �S�:�w߉�p߭ߔ���D�V�}����-�?�Q�c�u�)	��� ����������� ��� D�+�h�O�a������� ��������@R�9v	�`�Z��$U�I_POSTYP�E  `�?� 	 ����QUICKME/N  ����� RESTORE� 1 `�?  �i�!S`N�m~� �����/%/7/ I/[/�/�/�/�/�/ r�/�/�/j/3?E?W? i?{??�?�?�?�?�? �?�?O/OAOSOeO? rO�O�OO�O�O�O_ _�O=_O_a_s_�_(_ �_�_�_�_�_�O�_o "o�_Fooo�o�o�o�o Zo�o�o�o#�oG Yk}�:o��� 2���1�C��g� y���������d�����	��-��SCRE�� ?�uw1scHu2h�U3h�4h�5h�6h��7h�8h��USE�RJ�O�a�TI�j�k�sr�є4є5є6�є7є8ё� ND�O_CFG !����Ѩ PDAT�E ���?None _� ���_INFO 1"2`�]�0%3�x� 	�f�����˯ݯ��� ���7��[�m�P���ࣿ��ǿ�J�OFF�SET %� ԿσA֏�*�<�N� {�rτϱϨϺ�Ͼ� ���A�8�J�w�n� �ߒ�����
�����UFRAME � ʄ�G�RTOL_ABRT&��>�ENBG�8�G�RP 1&<?Cz  A���� ��������������:�� Ug��V�MSK  j�]�X�%N#���]�%�߫���VCCM�'����RG��*�	���ʄƉD � �BH)�p<2C�2)��PN?�` ��MR��20��p����"�р	 ���~?XC56 *�������N�5р��A@<C� ���ʈ)@;h�c���Rр|�Ђ B����6� t/T1/ /U/@/y/ d/�/�/�/�/*/�/	?��/???�c?u?��TCC��1��f�9��рр��GFSv�22w Й��2345678901�?�2ʈ"�6��?�!Oс>,12�QO_GB�@R 8N:�o=L����� ������OOA�O�O @O_dOvO�O�O�O�_ �O�O�___�_<_N_ `_r_Soeo�_Ro�o�_��_oo&o8o��4S�ELECF�j��$�VIRTSYNC� ��6�Bq�SIONTMOU4-tр��cu���3U��U��(�� FR:�\es\+�A\�o �� MC�v�LOG�   7UD1�vEX�с�' B@ ���qDES�KTOP-8U37T7F�6��q:�^��σ �  =�	 1- n?6  -��ʆ��xf,p�#�0=�̩ʹ���r�xTRAIN��2�1.���
. d��sq4w (,1��0�� )�;�M�_�q������� ��˟ݟ���I���crSTAT 5���@�o����E:$���ۯ�_GE��6nw�`. �
���. 2�HOMIN���7U��UC� �r�a�a�aCG��um�JMPER�R 28w
  ʯE:��suTs���� �߿���'�9�OϠ]ώρϓ�_v_�pR�E��9t���LEXr��:wA1-e��VMPHASE � RuCCb��OcFFLpc�<vP2�t�;4�04��8����b@�� �bb>?Gs33��Á�1�рL��ҕԈ�|��t�>x��Â�xf�o.���8/?P�X� $�2� x����0� ��� 6�+���l��\�j�|� ��������� �D� V���ZTf���� ������. �, BPb����� ��//(/:/� y/�b/��/�/L/ ? ??<?n/c?�/�/ �?�?�/�?6?�?�?�? OX?j?\O�?�OJO�? fO�O�O�O�O0O%_TO _xOm_�O�O�O�_�_ �_�__o>_P_EoWo �_xo�_�o�o�o�o���TD_FILTE:t�?�� ��Wp��]o$6HZl ~������ ��)�;�M�_�q�������SHIFTM�ENU 1@x�<��%����я�� 0���f�=�O���s� ����䟻�͟����P�'�	LIVE�/SNAPD�v�sfliv�b��{�ION G�yU���menu�����:�����±���A���	����b�K�S�5M����m`@�е���A�pB8��B����Ӝѝ�������m`� ;ӥ�/�M�E��uY��M�ֱ�MO��B���z���WAITDINEND�3���sOKN�.�OUT#�r�Sa�4�TIM�����GϮ�@π��`ϱ�ϱʞ�2�R?ELEASE���f�TM�����_ACTx��Ȫ�2��_DATA C��ի�%i��ߪ���R�DIS�b��$�XVR2�D��$�ZABC_GRPW 1E8�n`,@h�2��ǽZIP1�F�D� cCo������x�M�PCF_G 1G�8�n`0<o ���=�Hx8����t� 	�>w�  8R���0��e�����?�k�� ����5��
\�>�  �a � ����7������I��z��YLINuD�aJ�� �f ,(  *s��K�p���� �//+.mN/� r/Y/k/�/��/�/�/ 3/?�/�/J?1?n?U?`�/�?�?v�C�2K8��� ��O`o��7O~[Ol�?�Og���AA�ASPHE_RE 2LS�? �OX?�O__>_�?�O t_�_?�_I_/_�_�_ o�_]_:oLo�_�_�o �_�o�o�o�o#o l$7�ZZ� �k�