��   u��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����UI_CONF�IG_T  �� A$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]2�ODE�
3CWFOCA �4C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"��%�!BA�!j ?Ɵ"BG�%�!jIN=SR$IO}7�PM�X_PKT��"IHELP� M{ER�BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�; } &USTOM0� t $} R?T_SPID�,D�C4D*PAG� ?�^DEVICE�PISCREuEF���IGN�@$FLAG�@C�1 � h 	$PWD_ACCES� E �8��C�!~�%)$LABE� O$Tz j�@��3�B�	CUSR�VI 1  < �`�B*�B��APRI�m� t1RP�TRIP�"m�$�$CLA�@ ����sQ��R��R�hP\ SI�qW  �
�QIRTs1q_�P'2 �L3hL3!p�R	_ ,��?����R�P�S�S�Q��� , ��  o��
 ��zQQocouo�o�o�o�o Mo�o�o *<�o`r��� �I����&�8� J��n���������ȏ W�����"�4�F�Տ j�|�������ğ֟e� ����0�B�T��x� ��������үa������,�>�P�b��P_TPTX��򨸅����P sm����$/softp�art/genl�ink?help�=/md/tpm?enu.dgd��� �"�4��X�j�|ώ� �ϲ�A��������� 0߿�A�f�xߊߜ߮� ��O�������,�>�V���zQ'f	f�Sh�($�ߕ������������zQ�Q�op������v�Fc�n�(a��*������  ��P����@�v�n���8)��#`  �V������SB 1�XR_ \ }�%`REG V�ED�� wh�olemod.h�tm4	singl�Edoub\�triptbrows�@�! ����/A�S|�/Adev.sJl�o�1�	t���w �G/Y/k/5/�/�/�/8�/�/ ?� �P? *?<?N?`?r?�?�?�? �?�6�@?�?�?�? O 2ODOE	�/�/wO�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_ �_��_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	-?? z������� 
��O@�R�!�3��� ��QOcOI�ݏ�� *�%�7�I�r�m���� ����ǟٟ�����_ /�)�W�i�{������� ïկ�����/�A� S�e�w�����iֿ� ����0�B�T�f�x� s��Ϯ�}Ϗ����ϭ� ����>�9�K�]߆߁� �ߥ����������� #�5�^�Y�k�9���� ������������1� C�U�g�y��������� ������ſ2DVh z�������� 
��@R	�� �������/ */%/7/I/r/m//�/ �/�/�/���/�/?!? 3?E?W?i?{?�?�?�? �?�?�?�?OO/OAO SO!�O�O�O�O�O�O �O__0_+T_f_5_�G_�_�_�Z�$UI�_TOPMENU� 1�P�QR 
d�Q�fA)*defa�ultqOZM*�level0 *\K	 o� So��_Qocbtpio�[23]�(tpst[1�heo�ouo�3oEo�-
h58E?01.gif�(?	menu5&yp�Hq13&zGr%zEt4M{4�a����� ����eB�C�U��g�y�����,�pr�im=Hqpage,1422,1�� ݏ���%�0�I�[��m������2���c?lass,5��០���)�4���130�f�x�������5���53ʏ����( �2�5���8ٯm� �������4�ٿ����!�3�^I�P�Q�_ k�m]��a[ϕ�o�f�ty�m�o�amf[�0�o��	��c[1364�g.�59�h�a����tC8$|Gr2 uK}��azmWw%{�� �sK�]�6�H�Z�l�~� ɿ����������𢡊��80$�?�Q�c�u�����̐2�������� ��	��ʟ?Qcu �(T�������Ѥ1.�N`r������ainedic����/�/��confi�g=single}&��wintpĀ  /`/r/�/�/]J�QV� �/�/e�/�o�o?? 1?D?U?g?y?�?�/�? �?�?�?�?	OO-O?O �aO�O�O�O�O�O�O ��__*_<_N_`_�O �_�_�_�_�_�_m_�_ o&o8oJo\ono�_�o �o�o�o�o�o{o" 4FXj�o|�� ������0�B� T�f�x��������ҏ���MNS�,�wω� �����w���s��<����ϡ�u�͔�V�|�F7��7����԰�Οhp��ߔ�6��u7�� � �����/�A��227쯃������� ˿Z�l�����,�>�P�/!$13�ϛ� �Ͽ��ϐ�����+� =�O���s߅ߗߩ߻� ����"���'�9�K�]�����6d����0����,$۬74r�� /�A�S�e��,����%�	TPTX[2019�����24����������18������P�
����0P2��`�1_��E�tv��p���Q�u10��1=�ïqC:4$tr?eeviewA#��3�&dual=�oU81,26,4����n��� �	//-/�Q/c/u/��/�/�/ֺ;@b�3 `r�?)?;?F/_? q?�?�?�?�?�/�/\	2�/t2��O1OCO�?��1�/E���O�O��O�6XO��edit�zO�O_._@_׹ ?���OCL_�_�_�_ ~��_�_G�o}o� CoUogoyo�o�o�o�o /o�o�o	-?Q duӥ����� ��I?2�D�V�h�z� �����ԏ���
� ���@�R�d�v����� )���П������� <�N�`�r�����%��� ̯ޯ���&���J� \�n�������3�ȿڿ ����"��_�_X�o |��o��ϱ������� ���ߋ�)�S�e�x� �ߛ߭߿��ߓ�� ,�>�P�b�t￿��� ����������(�:� L�^�p���������� ���� ��$6HZ l~����� �� 2DVhz ������
/ �./@/R/d/v/�/7� IϾ/m��/I���?? )?;?M?`?q?�?�/�? �?�?�?�?OO%O7O ��nO�O�O�O�O�O�O %/�O_"_4_F_X_�O |_�_�_�_�_�_e_�_ oo0oBoTofo�_�o �o�o�o�o�oso ,>Pb�o��� ������(�:� L�^�p��������ʏ ܏/�/$��/H��? MOk�}�������ş؟ �W����1�C�U�h� y�����_Oԯ���
� �.�y�@�d�v����� ����M������*� <�˿`�rτϖϨϺ� I�������&�8�J� ��n߀ߒߤ߶���W� �����"�4�F���X� |��������e�����0�B�T����*default�a�2�*level8���������{�� tpst[�1]��yt?pio[23���u������	�menu7.gi5f�
�13�	��5�
��
�4�u6�
ʯ?Qcu� ������// �;/M/_/q/�/�/�/~6"prim=��page,74,1�/�/�/??+?6"��&class,130?f?x?�?�?�?=?O25�?�?�?O O2O5#D<�?lO~O�O0�O�O�/�"18�/�O@__'_9_DON26@_�u_�_�_�_�_��$�UI_USERV?IEW 1���R 
���_>��_
o�m(oQocouo�o�o<o �o�o�o�o�o); M_qo~�� ����%��I�[� m������F�Ǐُ� �����.�@���{� ������ßf����� �/�ҟS�e�w����� F�P���̯>���+� =�O�a���������� Ϳp����'�9�� F�X�j�ܿ�Ϸ����� �ϐ��#�5�G�Y�k� ߏߡ߳����߂��� ���z�C�U�g�y�� .������������ -�?�Q�c������� �������)�� M_q��8�� ���� 2� m���X�� �/!/3/�W/i/{/ �/�/J�/�/�/B/? ?/?A?S?�/w?�?�? �?�?b?�?�?OO+O �/�?JO\O�?�O�O�O �O�O�O�O_'_9_K_ ]_ _�_�_�_�_�_lX