��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  % � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d PPINFwOEQ/ ��L A �!�%/� H� �&�)EQUIP 2� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CES0s!_81F3K2> ��! � $�SOFT�T_I�Dk2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5Xk2S�CREEN_(4n_2SIGE0_?|q;�0PK_FI� �	$THKY�GPANE�4 ~� DUMMY1d�DDd!OE4LA!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTc@�D5�F6�F7�F8�F9�G0�G�GJA �E�GbA�E�G1�G ԂF�G1�G2�B��ASBN_CF�>"
 8F CNV�_J� ; �"�!_C�MNT�$FL�AGS]�CHE�C�8 � ELLSETUP � o$HO30IO�0�� %�SMACR=O�RREPR�X� D+�0��R{�T �UTOBACKU~�0 �)�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?��P�1E��#sAsTB�d��MO� ��cE D [Mp�c��^qREV�gBILrw!XI� ~QrR  � �OD�P�q$NO^PM�Wp�t�r/"�w� �u�q�r�0D`S p{ E RD_E�p~Cq$FSSBn&�$CHKBD_S�E^eAG G�"?$SLOT_��2$=�� V�d�%��3� a_EDIm  ? � �"���PS�`(4%$EyP�1�1$OP�0r�2�a�p_OK�;UST1P_C� ���d��U �PLACI�4!�Q�4�( raC�OMM� ,0$D ����0�`��EOWBn�IGALLOW�G (K�"(2�0VARa��@�2ao��L�0OUy� ,�Kvay��PS�`�0M�_O]����C�F�t X� GR�P0��M=qNFL�I�ܓ�0UIRE��$g"� SWIT{CHړAX_N�P]Ss"CF_�G�� �� WARN�M�`#!�!�qPLI��I�NST� CO�R-0bFLTR^C�TRAT�PTE�>� $ACC1a��N ��r$ORIأo"��RT�P_S�Fg CHG�0I���rTא�1�I���T�I1��� x i#�Q��HDRBJ; C,�U2'�3'�4'�5'�U6'�7'�8'�9{5;CO`T <F П�����#92��LLE�Cy�"MULTI�b�"N��1�!���0�T_}R  4F STY�"�R`�=l�)2`�����`T |� �&$c�Z`d�pb��P�MO�0��TTOӰ�Ew�EXT����ÁB���"�2� ��[0]�}R���b�}� D"}����Q0���Q�kc��A�^ȇ1��ÂM���P�� ŋ� L�  ���P�z�`A��$JOBn�x/�i�G�TRIG�  d�p�߻��� ��7�����'��_�M�b! t�pF̝ CNG AiBA � ����M���!���p � �q��0��P[`��,i�*�"6���0t�B񉠎"J��_Rz�gC�J��$�?�Jk�D�%C_�;������0ФR�t#�C ������G����0NHANC̳$LGa��B^a��� �D��A�`��gzRɡ�!��p�3DB�RA�sAZ�0KELT��\���PFCT&��1F�0�P��SM��cI��1�% ��% ��@R��a���� S��&���M 00{o Ve#HK~�A^S��h�����I_T$�"�6SW�CSXC�)�?!%��p)3��T�$@��PANN�&�AIMG_HE�IGHCr�WIDLI AVT�0��H F_ASPװ��`�EXP�1���CWUST�U��&��
|E\�%�C1NV q_�`�a��' \%1y�`OR�c,"�0gsdk��PO��LBSYI�G��aR%�`좔Psp�m��0k� PXW�ORK��(~!$S�KP_�`maJ0D�B<qTRp ) ���P���� �0f�DJ!d/�_CN�0�R�#� �'PL�S�Q��d�s�DKA7WA�w'�^A�@NFZp ML�DBU��*�"&!PRS�7�
ЖQ�����+ [pr��$1�$ZϢ�LBi9,v?�3ʠ��-�?ʮ4C��.�?�4EN9Ey��� /�?�3�J0RE`��20Hz��CuR+$L,C�,$i3
�? =KIN�E@�K!_D�I�RO�`����ȳqvC���h �FPAÃ3uRf�PRN�B�MR���U!�u�CR[@EWyM �SIGN���A� .q�E�Q-{$P��.$Pp &2�/ P7�PT2�PDu`L���VDBA|R@�GO_AW����Jp � �DC�S�pZ�CY_ �1���@1<�Q?fI+G2�Z2>fN>������
�qS&c}P2 P7 $��RB?�e�eP=hPwg�QBYl��`gT+1�THNDEG�23��KS�SE|�Q��SBL�Y�cc�T�qrRL�4 �HpZ ���VTOFB�l�FEfA�ǿbh�TqSW5�bDOC���MCS�f�`Z$(r�b H� W0��T�K�rRSLAV�16�rINP��f���LyqQP�7� $,�S���=��v�,�uFI��r� �sc�!��!W1ԭr'NTV'��rV	��u7SKIvTE�@W0���:�J_� y_�00�SAFE��A�_SV��EXCSLU��B �PDJ 	L1�k�Y�d�ƻr�I_V� !PPL1Y 0b���DE~w���_ML2�B $VORFY_�#��Mk�IOU��憻 0���2:�O�P��LS�@jbF;�3572��Sr�� Px%X�{P�hs� Ή� 8 @� TAx� qঠ �c/_SGN��96��� �@�A�����iPt!0��s"��~UN�0jd Ք�U���B �@�  ��� ����!l�wOGI�2: @�`1Fؒ���OT�@@Ð:41(�77471�M`NI�2;�R����r��A�q��DAY1#LOAD�T/4~�;3�0� �EF�XIJ�b< @%1O�|�3� _RTRQ��G= D�`@��Q@  �EjP"�㥂��<�B�� 	�@��GAMP��]>��a�����a�8Sq�DUt�@q���"CAB���?A��0NSs���IDI�WRK�^�� �V�WV_]���> ��DI��q�@�� /.�L_SE2�T���/�Z`��0��#�E_��u�v�j��SWJ�j� 𐲰��	���=c�O�H�z�PPJ�v�I	R!��B� ��w�d�p�B"����BASh���� X ���V����?�C��Q��RQDWf��MS���AX}�<8�u�LIFE� �7�A1C�NJ���S��DH���Cs�>��C`QN"�U��3OV� _�HE����'SUP�hbC�� _�Ԥ���_����[Q
��Z��W���ו�Tb��XZ$ `1��+Y2F�CM@T��t@r�N�p���;CT9A `�P.�sHE��SIZy���u��BN�pUFFI���p� �Q/4�0�<26711�MS�W9B 8�KE�YIMAG�CTM�@A��A�Jr�>1�OCVIET���'C ��V L�t����s?� b� :D��"pST�! x�0�� 0��Ѡ��0�>��EMAIL���@�����c`_FAUL⍢EH�CCOU��p}!��T@��FO< $���eS]�v��ITvBUF�砤q���T  ���BdC�t����#��SAVb$)�e�A� }���Pi�e@�U�b`_ H���	OT{BH�lcPր(0�
{��AX1#�� �@��_GJ�f1YN)_�� Gj�D�U/0�e��M����T
8�F��ِ�A!�H�(@u���C	_r@�@K�D�����=pR���uDS�P �uPC�IM@b��J���U�0�ЁEƀ��IP�sun��D  �TH0ȸc��TuA�HS{DI�ABSC�ts��0Vzp*} �$,�#��NVW�G�#�$H0� FJ�/d�j�ASC��U��MER��uFBC3MP��tETH�!AmI��FU��DU 0�a�@;⠂CD�O �� ���R_NOA�UTg` J�`�Pp2��n4ĥPSm5�CF }5CI�.���k3� =KH *}1Lp��Q��& �I���4#Q�6s��6@ѡ�60��6���67�9�8�99�:J��8�:1�J1J1J1+J1�8J1EJ1RJ1_J2RmJ2�;J2J2JU2+J28J2EJ2RJU2_J3mJ3�:3KBJ3J/�G8J3EJ�3RJ3_J4mB|�ESXT�>aLC`���F�fF�5Q9g�5�3pFDR�MT��VC��C�wa}".C�REM,�FAj�OVM��eA�iT7ROV�iDTm �jMX�lIN�i���jN�IND�`!�
x<p /$DG�Ð�`opS�9�D��`R�IV)0Qbj�GEA-R�IO0�K�bu�Nj�x�.؎��p�q>j�Z_MCM>�C��d`��UR)2N ,<{1��? ��
 s?�pI�?�q	E���q%1�T0lb�Oߠ��P� �R�IT5��UP2_� P Ѡ#TD = ��C����qP�J�0��$BAC;Q TЕ�$9 O�)��OG�%E��3e&0IF�I��e0�0����PuT��MR2ie�R vbY�vbLIq��{g�����f��Ŗb_mADN~F�_F�I4+�M;v|`r}DGCLF��oDGDY��LD�q�>t5[�5S�كk�S���M� T�F9S� l�T P�)����
�/$EX_)�@�)�1�� ��*�53b�5b��G�!iegU � p&2SWK}O��DEBUG�SL��0�GRY�zU�#�BKU� O1�@ O�PO8��Π�0��ΠMS]�OO,��SM]�Eq�1�pQ`_E V �$�X�c`TERM�2�W;�ype�O�RIĀ6�X;�4&�SM_��$7��Yk�TAy�Zk�U}PB�[� -���QbV$G���W$�SEGźאELT}O��$USE0NFI����p����`���X$UFR�����q0豈�D5h�OT1Ǵ TA_ �C�wNSTd�PATT!<��Y�PTHJ!B0�En�K0�ART�� ��������REyL��&SHFTF"��_���_SH��M��!B0x� ��n���Z����OVR
#&SSHI����U�2 ��AYLO$ 5I�1�_�d���d�ERV�0*�} ��b?�d���Q����A��RC<
���ASYMh��F�WJ�apE�����f�2�U��d�5����D5��P#Gи!�	�ORd�M���!���\��΢�^���D���k�] �tE���TOC�1졳q��OP��N Pz�3&1���aO�a�> RE��R�#&OX0��`�e��R]���������e$PW�RSpIM��[�R_���VISy�r����UD����� �^>�$H����_�ADDR9fH$�G a�z�s�i1R� .=_ H8�S� ��S��C��C��CS)E�aY�SO0���` $���_D�`���PR��r�HTT� U�TH�a ({0O�BJE1u���$�9fLEP�-=b� � *g!AB%_qT��Sk�#�DBGLV5#KR�L"�HIT�BG�0LO���TE�M4$��b������S�S�p�4JQUER�Y_FLA��f W(YA���c��� 3PU�"B�IO0���4G��H��HB _�IOLN~�d/0�i�C��$SLz�� PUT_�$���Pwp�rwSLA�� e/2@����ӡ���0{IO F_AS�f��$L��U�� �#�04�#����,ЃHYOgN!'#�1 U;OP�g ` l!�9f�b>$�`E&�!��P�����'�!E&�"�&~�P_MEMBk0�T h X IPz�v��"_#0v�����0��Oc6�1w�D�SP�' $FOC�USBGv�D�UJhfi � 60S���JOG�W2DIS��J7��O��$+J8�97��I6!�2>�77_LABQ���x�0�8�1APHI�p�Q�3�7D+�J7�JRA4`P�_KEY�p �KIL�MON�j&`$�XR =0cWAT�CH_ �DӘ�U1E�L� �y�B�k� GpG�VP�-ffBC�TR��fB5��LG|�l ��+h�"��?LG_SIZ{Y�`�E
��F
 �FFD�HI�H�H��F�HM��F �@���C5V
�5V
 5V �@5VM�5W�`S)@S�H���@Nv1��mx � ��R��4a�PÀ�U�Qk�L�S�RDAU�UEA I���R�PGH���AO�GBOO~�n�3 C-"2�ITGcdܝ�)&REC-jSC�RN)&DI(#S��RG����cl� !#��b�!Sa"�Wkd!�T!#JGM��gMNCH"F�N�2�fK�gPRG��iUF�h	��hFW�D�hHL/ySTP��jV�hĀ�h`�hRESgyH!�{&C�@Es��!#���g�yU�t�g�¬f|@6#�bG�i4�PO�JzZeEs�M�w82�iEX'TKUI�eIP�cw� �c���c���`�a���`�s��Jg��KaNO{��ANA"貇�VA�I�0zCL����DCS_HI������b��O����SI)�r�S'��hIGN�@���C�aT����DEV�wLL�єQ6@SBU𠔠oa@�mT��$�GEM'P9nD,�EsAb�pa@�ЅC�!��OS1��2��3��)Ж�����q �T0v-�p絡.e�IDX����-fL�b�ST�m R�PY0���� _p$E��C���  ����� ��r L*</��Q(6����6�EN 6�Օ~Kc_ s Y���P$ dKaD� �M�C�Rt �T0C�LDPm ��TRQ�LI`��e0x�f�FAL>1��_����DUA���LD������ORGe0�r���WX������Y���V�O�u �� 	���uu���Si�Tx��00�ްS�}[�RCLMCi�����{�m[�ՐMI���O�v d�Q6�R�Q�00�DSTB���Y� ��{a��A�X��@�� �EXC+ES����M��w(��¹�a��j��x(��_A�ʠ� l����V�K|�y� \*�2��$MB�LIE��REQGUIR����O��ODEBU��L�M{�zW�.!��B��Di�+�N,03Ѩ�{�R��RkHV�DCE��TIqN3 `!�TRSMw0�p�S�N�����s<�P�ST�  |h�L�OC9�RI� 9�E�X��A��:�����O�DAQo%}��$@�Q΂MF�A��_���p�C��P��SkUP�
C0FX���IGG�"~ � 0��MQ���v�5@� %����m ��m ��<��6#DATA����AE� 1�NP" N��� t�MDI�F)?�!��H����1!� �Q"AN�SW�a!ܑS�!D��)��H3Q�$� -?�CU�@V_ >0L���LO�P$�=�$����L2�������RR2I5�O  ��QAX�� d$CALI���NUG�2gRsINp<$R�SW0��K�AB�C�D_J2SE�����_J3v
�p1SP�@6 ��P�p�3��\���B�J���P�O���IM��[�CSKP ��$�P�$J�Q[Q,6%%6%,'��_cAZW��h!EL��<���OCMP�����1X0RT�Q�#�11�c@�Y�1��(�0:�*Z�$SMG�p��L��ERJ�[IN� ACߒ���5�b��1�_B��542d�[�n�14X҆f>9DI~!��DH �t30���$Vlo�Y�$�a$�  ��A�<�.A�����H �$BE�Ly lH�ACCE�L?��8���0IR�C_R��R��AT<w�c�$PS �k�L�yP D��0Gx�Q�FPATH�9�WG�3WG3&B��#�_@�2�@�AV���C;@��0_MG|a$D�D�A@[b$FW�(����3�E�3�2�HD}E�KPPABN.GROTSPEE�B���_x�,!��DEF�g��1�$USE)_��Pz�C ����YP�0V� �YN���A{`uV�8uQM�OU�ANG�2�@O9LGC�TINC~����B�D���W���ENCS����A�2��@INk�I&Be���Z�, VE�P'b2�3_UI!<�9cLOWL3��pc x��UYfD�p��Y�� ��Ury�C$0 fMOS`�Ɛ�MO����V�PE�RCH  vcOV�$ �g9��c��\bYĀ���'�"_Ue@0��A&BuLcT����!epc�\jWvrfTRK�%h�AY�shчq&B��u�s���&l��Rx�MOM|���h�ﰞ �Ą�C�sYC���0D�U��BS_BCKLSH_C&B��P �f�`}S�7��RB��Q.%CLAL��b?�8�pX�t�CHKx�H��S�PRTY�����e�����_~��d_�UMl�ĉCу�ASsCLބ PLMT��_L�#��H�E ������E�H�`-��Q#p_��hPC�aB�hH��ЯEǅCw���XT�0�GCN_b(N�þ���SF�1�iV_RG�e�!�� r����CATΎSH ~�(�D�V��f�0'A�	� �@PA΄�R_Pͅ�s_y�뀎v`�`x��s����JG5��6Ф�G`OG���rTORQUQP��c�y��@�Ңb�q�@�_W �u�t�!�14��33��3�3�I;�II�I�3F��&������@VC"�00���©�1��2�8ÿ�¶�JRK�����綒 DBL_SMt�QO�Mm�_DL�1O�GRV:�3ĝ33��3�H_��Z@a��COSn˛ n�LN ���˲��ĝ0��� �� e��ʽ̃��Z���f��MY���z�TH|��.�THET0beNK23�3Xҗ3��[CB]�CB�3C��AS���e��ѝ3���]�SB�3��h�GT	S@! QC���'y�x�'����$DU�� ;w	��Q�����q9Q����$NE$T�!I�����)I7${0LсAP�y��`�k�k�LCPHn�W�1eW�S�� �������W���������{0V��V��0��UV��V��V��V��UV��V�V�H��@����7�����H��UH��H��H�H��O��O��OF	��O���O��O��O��O*��O�O��FW�}���	�����SPBA�LANCE�{�LmE��H_P�SP1��1��1��PFULC5\D\��:{1��!UTO_���ĥT1T2��22N���2, ����q^P<�-B#�qTHpO~ |�1$�INSEG�2�{aREV�{`aD3IFquC91�('o21�dpOB!d�=���w2��7P���LC�HWARR�2AB����u$MECH`��ДQ�!��AX�q�PB��&r�~2�� �
�"��1eROBF�`CR r�%��%x0�MSK_�4� WP �_OPR�1�2(47Qst1�,`*R`(0)cB�(0|!IN!��MTCOM_�C���0�  ��@0 �A$NOR�Ec�2�l ~2�� 4�GR��%F�LA!$XYZ�_DA��LP;@DE�BU�2 �0lR�0�u ($mQCODS�G �2�r� �p�$BUFIND�X*P0;@MOR3� H%0�p�0���:@�p�QB�"�1c��NF�TA9Q�#C�rG.B� �� $SIMU�L���0�As�AsO�BJE3�FADJ�US�H�@AY_It��xD�GOUTΠ��4�p�P_FI�Q=8AT#�Y,`W�1�P +�PQ+ 9�uDNjPFRI �PUT0��RO�
`E+�Sp��OPWO��0�},@SYSBUi� @$SOP�QBy��ZU�[+ PRUN,n2�UPA;0D�V�"��Q�`_�@F��PP!A�B�!H��@IMAG�S�%0?�P!IM�QAdIN$��RcRGOVRDEQ�R�@��QP�Pc�� L_`��feÂސRBߐ�<pX�MC_EDT'@�  H�Ni M�b<G��MY19F�0�EaSL30� x $OVSL�wSDIsPDEXǓ��f֓Hq�bV+��eN �a
��Pp�cwx�bzw��d_SET�0� @�Cr�%9�SRI�A3�
Vv_��bw{qnqf��-!�@� �4BT� àA�TUS�$TR�CA�@PB�sBTM$�w�qI�Q�d4F��s\�`0� D%0E�P�b�rr�E1"�qQpd��qEXE�p���a�"��tKs�Rp&0�p3UP�01�$Q `XNN�w���d���y� �PG|5�? $SUB�q�%�xq�q|sJMPWAeI$�Ps��LO ���1
 �E$RCV?FAIL_C@1�PÁR%P�0�#���Ȕx� �
�R_PL|s�DBTBá���PB3WD��0UM���IG�Q `�,�TNL ��b�ReQ�2��$�qP��@EǓ��|֒��DEFSP� � L%0� ��q_���CƓUNI�S��wĐe�R)��+�_uL
 P�q���H_PK�5��2RETRIE|s�2�R�"@���FI�2� Ϙ $�@� �2��0DBGLV~�LOGSIZ�CH� ���U�"|�D?��g�_T:��!M�@C,
 #EM��R��y0>�8CHECKS�BS�Po01��0.��0R!LbNMKET(��@�3�PV�1�� h�`ARp� ��1)P�2>�S�@OR~|sFORMAT��L�CO�`q����$�Z��UX�P!r?qP�LIG�1�  ˣSWIm �a|A���,�G�AL_ G� $`@��B�a��CS2D�Q$E�1��J3DƸ�{ T�`PDCK�`|�!LbCO_J3�����T1׿� ��˰C_Q�` �; ��PAY��S2�u�_1|�2|�ȰJ�3�ИˈŬƗ�tQTWIA4��5��6S2MOMK@��������4��y0B׀AD���������PU��NR���C���C���4�` I$PIN� u�41�žӁ�:q�R ~ȇ��ٯ��:�h��a�֬��ց�1�'1R�\uSPEED G ��0�؅��7浔؅� %P7�m�F��U��؅SAM =G��7��N؅MOV	B� e0 �� ��c2��v��浐 �� ���c2nPsR����dİ$QH���IN8� İ��?�[�6�؂A���xX����GAMM|�q�4$GET1R�@�SDe�mB
�L�IBR[�y�I�7$HI�0_5a@c2�E`@#A@ 1LW^U@	�1a��&o�ʱC=�n S`�po �I_�� pPmDòv�ñ'�����mD��	ȳ ��$�� 1��0I
zpR� DT#|"c���~ LE^141�qwa��?�|�MSWFL��MȰSCRk�7 �0��Ѻv���Z 0�P�@9@����2�cS_SAVEc_Dkd%]�NOe�C�q^�f� ��uϟ� }ɕQ��}���}*m+��9��ժ(��D�@���� �������b31�RA�Mam�7
5�#��^����Mtա � F�YL��
A'�VAS	BtRna`7GP�B
B�l3
A%`�GSB1W? �2�2cЬ3oBB1M&@�;CL�8���G$�b�1v���M!LrǢ �N�X0�d$W @�ej@b�� @=� BD�BK�B�-�> @�P����ycİX �	OL�ñZ�E���uԷ� ��OM �R/d/v/�/�/��A�XjM`�aPLe�_��� |��H ��jV ��yV��yP�ʗW�V��9E��� IW���8���NTP=���PMpQU�� �� 8TpQCOU�,�QTHQ�HO�Y2`HYSa�ES���aUE `"#�O.���   �P�0��rUN�p�3��O$�J0� P�p^e��x����OGRA�q�k22�O�d^eITxm�aB`INFOI1����k�ak2��O�I�b� (!SLEQ(��a��`�foayS� ��� 4Tp�ENABLBbpPTION|s����Yw���1sGCF��O�c$J�ñfb���R�x!�]ot �QO�S_EDŀJ0� I�N��@K�᪃�ES NU�w�xAUyT,!�uCOPY��P���v�8 MN����PRUT�� ��N�pOU��$�Gcbn�l�RGAD5JI1�2�X_B0ݒC$ ����@��W���P�����@㊀��E�X�YCLB��N�S6u�N0�LGO��A�NYQ_FREQZ�W���+�p�\cLAm"����Ì��uCRE  c� I�F�ѝcNA��%�i�_GmSTAT�UQPmMAIL �� 1��yd����!���ELEM�� ��7 DxFEASI Gq2��v��q!�er$�  I�`�"��0ae�|I�ABUq��E�`D�V֑a�BA!S��b� [�Ub�r �% $y���RMS_TRC�ñj�� �Ca��ϑ��,r���C��YP	 � 2� g�DU���� �Ԣ�0-�1��1���NqDOU�ceNrs���PR30;p�rG�RID�aUsBAR�S(�TYHs�a#�O\�I1� Oa_���!ƀ��l�O�@7t�� � �`�@PO�R�cճ��ֲSRV���)���DI. T����!��+��+�4�)�5)�6)�7)�8���QF��:q�M`$VALU|�%��ޡ��7t�� Cu'!�a���� (gp#AN#��R�p0�> 1TOTAL��[і�PW�It�&�R�EGEN$�9��SX���sc0��Q���PTR��Z�$�_S ��9Ђ�sV���t���rb�E���x�a�"^b�p��V_H��DA�C����GS_Y4!�B<�S�{AR�@2� f�IG_SEc���2˕_b`��C_�����w��?r��%�b�H�SSLG#�I1��p" =���4��S�2̔DE�U!Tf.p���TE�@���� !a����Jv�,"��IL_MK��z���@TQ�P�a���*�2VF�CT�P����^�Mu�V1t�V1���2��2��3��3
��4��4����С`���1�"IN	VIB@N�; �!BU2>2J3>3J4>4JI05���"�p�MC_YF`3 � L!(!�r�M= I��FM� [PR�� �KEEP_HNA�DD�!f�C�A��!����"O�Q I����"��\?�"REM9!��ϲ^uzU��e�!HPWD  }SBMSK�G�a	!B2B�
#COLLAB�!���2�����o��`I�T��A`��D� �,pFLI@��$�SYN� ;,M�@C�>��%�UP_DL�YI1�MbDELAhm ј�Y�PAD�A��PQSKIPNE5� ��``On@cNT�1� P_`` �b�'�`�B]0�'���) 3��)��)O��*\��*@i��*v��*���*9O�J2R‎��?sEX��T%�|1�{2�ܐ�|1�a��PRD]C!F� ��pR�sR�PM�'R^��:b�2�RGE�p2��3d�FLG�Q�J�t��SPC�c�UM_||0��2TH2NP��F@o0 1� m�0EF�p11��� l[P�E-Ds#ATWo�[�w�B�`��d�A�p3�BfcAHPnP�B��_D2gB�mO@O�O�O�O�O�G3gB��O�O_ _2_D_�G4gB�g_y_�_�_�_�_�G5gB��_�_oPo,o>o�G6gB�ao@so�o�o�o�o�G7gB��o�o&8�G8gB�[m�����ES����\@@ǡ`CN�@�!uE��^� @o��m�IO�ፉI��Ы2��@WE!� �W�: �1���0� y�5%Ȃ$DSB;���֒ �h CL@�­0�S232s�� ��0�u.��ICE�U{���PEV@��P�ARIT�њ�OPyB ��FLOW��TR2�҆]���C�UN�M�UXTA����INTERF�AC3�fU���	�CH�� t`� � ˠE�A$��&��OM��A�0נ�I���/�A�TN���Tо ��ߓ��EFA� �"!�Ґ�G� u!��� O��� &*�� ������  2� ��S�0�`�	� �$3@}%:B�Ŏ�r�_���DSP���JOG��V�h�_P�!s�ONq0%�0�z��K��_MIR����w�MT7��AP@)�w�>@"���;AS�������;APG7�BR�KH����G �µ! ^���i���P��Ҏ����BSOC��wNl���16�SVG�DE_OP%�FS�PD_OVR�du �DвӣOR޷�pN��߶F_�����OV��SF�<���
�F0����UFR�AF�TOd�LCHk"%�OVϴ ��W[ ���8�Ң�͠�;�  @ BTI�N����$OFS2��CK��WD����`�����r���TR�9�T�_FD� �OMB_C �B���B����(�.Ѻ�S�Ve��琄�}#�Gl)�<�AM��B_��jթ�_M@�~���<����T$CA����uDe���HBK�,����IO��թ���PPA���������Տթ���DVC_DB��?����A��@,�X� b��X�3`�@���3�0����ϱU�����CAB�0��ˠ���c� �Ow�UX~��SUBCPU�ˠS�0�0�R����!��A�R�ł�!$HW_Cg@A��!��F���!�p� � �$U� r�l�e�ATT�RI��y�ˠCYC�����CA���FLT ��������A�LP׫CHK�_�SCT��F_e�F1_o����FS�J�j�CHA�1��9I�s�8RSD_!聂��恩�_Tg�7��L �i�EM,��0Mf�T&� @�&�#��DIAG��RAI'LACN���M�0� "��1���L��{�kPRB�S   �p�C4�&�	��FU�NC�"��RIN��0 "$�7h�� S	_��(@��`�0��8`A��CBL� uA����DA`p�a���LDܐ ð�����j���TI%��@�$?CE_RIAA��+AF�P=�>#��D%T2� C��a�;��OIp��DF_L�c�X��@�LML�F}A��HRDYO���RG�HZ 7��|��%MULSE� p�����k$Jۺ�J����FAN_�ALMLV�1W{RN5HARDr���Fk2$SHADOW|�A���O2sƐ0N�r�J�_}���A�U- R+�TO_SBR���3���:e��6�?�3MPINF�@{��4��3RE�G�N1DG�6CV���s
�FLW��>m�DAL_N�:�@����C	����a�U�;$�$Y_Bґ� u�_�z��� �/�EGe���ðF�AAR������2�G�<�AXE��R�OB��RED��W�R��c�_�M��SY�`��Ae�VSWWR1I���FE�STՀ��(��d��Eg�)��D-�{2��BUP��\V���D��OTO�1)���ARY���R����6�נFIE����$LINK�!GT5H�R�T_RS��q�E��QXYZ�:�Z5�VOFF���R1�R�X�OB��,�8d����9cFI@��Rg��􃻴,��_J$�F�貿S��q0kTu[6��1�w �a�"2�bCԀ+�DU�¤F]7�TUR0X#��e�Q�2X$P�ЩgFL�Pd���@p�UXZy8���� 1�)�%KʠM��F9��8�ӓORQ���LfZW30�B�OP�d�,��t����A�tOVE�q_BM���q^C �udC�ujB�v�wL�wg��tAN=�Q�q D!`A�q��=�}��q�u��q���dC��"���E)Rϡj	�E��T�$ńAs�@�UeX`��W����AX�� F����N�R��+� �!+�� *�`*��`*�@�`*�Rp*�xp*�1�p *�� '�� 7�� G��  W�� g�� w�� ��� ���� ��đ��DEBU=�$8D3�h����RAB������s9V��<� 
��i� `A��-񷧴������ a���a���a��Rq���xqJ$�`D"�R9cLA�BOb�u9�F�GR�O��b=<��B_ ���AT�I`�0`���p�u���1��ANDfp��ຄ���U���1ٷ  ���0�Q������P�NT$0M�SERsVE�y@� $%`�dAu�!9�PO ��[0ЍP@�o@*�c��x@�  $.]�TRQ�2
\��B2f��j�D"2�{�" ~� _ � l"�T�c6ERRub�I���VO`Z���TOQY�V�L�@)�1R�Ƅ %G;�%�Q�2 [�T0�e�� ,7�ř���]�RA#� 2֓ d@����r� �Y@$�p�t ���OC�f�� � ��COUN�TUQ�FZN_C;FGe�� 4B�F��Tf4;�~�\� �
�xӭ�uC� ���M: �"`A��U��q: ��FA1 d�?&�X��@=����_B�A<�����AP��o@HEL�@��� 5��`B_BAS�3RSSRF �CSg�!��1
ש�2��3���4��5��6��7r��8
ל�ROO��йP�PNLdA�cAqBH�� ��ACK���INn�T��GB$Upq0� +\�_PU��,@0��OUJ�PHH����, u��TPF?WD_KAR��@&��REGĨ P�P�n]QUEJRO�p�`2r>0o1I0������P����6�QSEMг�O��� A�ST�Yk�SO: �4DI�w�E���r!_T}M7CMANRQ���PEND�t$K�EYSWITCH����� HE�`BoEATMW3PE�@CLE��]|� U���F>��S�DO_�HOMB O>�_�EF��PR>a9B�ABP�x�CO�!��#�O�V_M�b[0# IOcCM�d'eQ�v��HKxA� D�Q$G��Ue2M�����cFORCCWcAR�"�Ҋ�OM�@ � @r�:#�0UUHSP�@1&2&&E3&&4�A��s�O���L"�,�HUNLiO��c4j$EDt1�  �SNPXw_AS��� 0+@� @��W1$SIZ��1$VA���M_ULTIPL��#�! A!� � �$��� NS`�BS��ӂAC���&FRI	F�n�S��)R� {NF�ODBU$P ���%B3=9G�Ѫ�ny@� x��SI���TE3s�r�cSGL�1T�R$p&�П3a�<P�0STMT1q�3�P�@5VBW�p�4S�HOW�5��SV���_G��� Rp$�PCi�oз��FBZ�PHSP' Av��Eo@VD�0vC�w� ���A00޴ RB% ZG/ ZG9 ZGC �ZG5XI6XI7XI8*XI9XIAXIBXI  ZG3�[F8PZGFXH��TXdI1qI1~I1�IU1�I1�I1�I1�IU1�I1�I1�I1�IU1 Y1Y1Y2WIU2dI2qI2~I2�I2�I�`�X�IQp�X�IU2�I2�I2�I2 Y�2Y2Y�p�hdI3�qI3~I3�I3�I3��I3�I3�I3�I3��I3�I3�I3 Y3�Y3Y4WI4dI4�qI4~I4�I4�I4��I4�I4�I4�I4��I4�I4�I4 Y4�Y4Y5�y5dI5�qI5~I5�I5�I5��I5�I5�I5�I5��I5�I5�I5 Y5�Y5Y6�y6dI6�qI6~I6�I6�I6��I6�I6�I6�I6��I6�I6�I6 Y6�Y6Y7�y7dI7�qI7~I7�I7�I7��I7�I7�I7�I7��I7�I7�I7 Y7�Y7T��0Pz� Uc�� l�Dנ��
>A820��5��RCM2����MT�R��|���Q_��R-��ń����[��YSL�1�� � �%^2��-4�'4�-Y�BVALU��Ձ���)���FJ�IgD_L���HI��9I��LE_���f��$OE�SAbѿ� h 7�V?E_BLCK�|�1'�D_CPU7� � 7ɝ �����E����R � � �PW��>�E ��LA�1Saѝî���RUN_FLG�� ������� �����������H���Ч�|�T�BC2��� � _ B��� br� 8W?�eTDC�����X��3f�S�TH�e�����R>�k�ESERVEX��e®�3�2 �d��� ��X -$��L�ENX��e�Ѕ�RyA��3�LOW_7��d�1��Ҵ2 �MO$/�s%S80t�I��"�`ޱH����]�DEm�41LACE�2�CqCr#"�_MA� pl��|��TCV����|�T�������0B k�)A�|�)AJ��%E�M7���J��B@k�X�|���2p �0:@�q�j�x JK��VK�X�����ы�J0l����JJ��JJ��AAL���������e4��5�Ӵ N1��P ����LF�_�1�� �CF�"� =`�GROU���1��AN6�C�#\ R�EQUIR��4E�BU�#��8�$Tm�2���|ё �%�� \�APP�R� CA�
$O�PEN�CLOSD<�Sv��	k�
�.�&� �<�MhЫ�8��v"/_MG�9�CD@�C ��DB{RKBNOLDB>�0RTMO_7ӈ$r3J��P��� ������������6��1�@ �|�$��� �� ���'��-#PATH)'B!8#B!�>#�� � �@�1SCA����8IN��U�CL�]1� C2@UM�(Y"��#�"�����*���*��� PAYL�OA�J2LڠR'_AN`�3L��9�
1�)1CR_F2gLSHi2D4LO4��!H7�#V7�#ACRL_�%�0�'�$��9H���$HC�2�FLEX��J#�� P�4�F߭�����0��� :����|�HG_D����0|���'�F1_A�E �G6�H�Z�l�~���BE����������� �*��X�T,�C���@@�XK�]�o�^Av�T&g�QX>�?��4TX�� �eoX������������ ������	-	Ҡ�0@� �/�M_q�~�۠AT�F�6�E�LHP���s�J� �v� JEoCTR�!��ATN���v|HA_ND_VB��1ܟ�$� $:`F24Cx���SW5�� $$M,0 0�_Y�ni��P\����A��� 3�����<AM��_AmA�|��NP�_DmD�|P\ G��E�ST�aM�nM�NDY ��� C����0��>7 _A>7Y1�'��d�@i`�P��������""J$�� �O�4D'"��J���A'SYMl%A�� l&!��@�-Y1�/_�}8 � �$��� ��/�/�/�/3J	<�:;�1�\:9�D_VI�x�|��V_UNI�����cF1J����䕶� Y<��p5Ǵ�y=6��9 ��?�?>�wc�4�3�  �$� AS�S  ����s�  ��{�h�VE�RSIONp��~��
��IR�TU<�qσ�AAV�M_WRK 2 ��� 0  �5z��������� ��	8�)�L�{����:�w�^�|�(ܛݧ��7ѭ���������BSwPOS� 1��� <�� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������//�1/C/U/ⰑAXL�MT��X#�%�  dj$INs/�!i$PRE_EXE�(A� �&)0�q��������LARMRECOV �ɥ"
�LMDG �����[/LM_IF �ˆ!X/c?u? �?�?�:Q?�?�?�? OM, 
0�8O�4��cOuO�O�O�NG?TOL  ��ЏA   �O�K��P�P)�O ;� ?6_,_>_P_{� $BR_�_w�o_�_�_ �_�_�_o�_'oo7o]o�!��O�o�o�o�o �o�o�o+=O�a�PPLICA�T��?��� ��%@Hand�lingTool� �u 
V8.?30P/33�@lt���
883�40�slu
�
F0�q�z{�
�2026�tlu���_�7gDC3�pJ  �s�Nonelx� �FRA�������B�TIV�%�s�#��UTO�MOD� E�)P�_CHGAPON������ҀOUPL�ED 1��� ���"�4�uz_CUREQ 1��S  � >�>�*����4��!��x��~� ��u���Hm����HTTHKY����w���7� ���%�C�I�[�m�� ������ǯٯ3���� !�?�E�W�i�{����� ��ÿտ/�����;� A�S�e�wωϛϭϿ� ��+�����7�=�O� a�s߅ߗߩ߻���'� ����3�9�K�]�o� �������#����� �/�5�G�Y�k�}��� ����������+ 1CUgy��� ���	'-? Qcu����/ ��/#/)/;/M/_/ q/�/�/�/�/?�/�/ ??%?7?I?[?m??���P�TO�@����DO_CLEAN܏|��CNM  �K >�aOsO�O�O��OD�DSPDRY�RO̅HI��=M@ NO_'_9_K_]_o_�_��_�_�_�_�_�_J�MAX�p�4�1���a�X�4"��"���PL�UGG���7���P�RC�@B;@?K�_�_ebOjb�O��SEGFӀK�o�g�a ;OMO'9K]�o�aLAP�O~Ǔ� ������/�A��S�e�w���΃TOT�AL-fVi΃USE+NU�`�� ������P�RGDISPWMMC�`{qC�a&a@@}r��O�@f��e��_STRI�NG 1	ˋ
��MĀS���
`�_ITEM1j�  n�������� ��Ο�����(�:� L�^�p���������ʯ�ܯI/O S�IGNALd��Tryout M�odek�Inp��Simulat{edo�Out.�OVERR�@� = 100n�In cycl"��o�Prog A�bor8�o��S�tatusm�	H�eartbeat�i�MH Fauyl����Aler�� �ݿ���%�7�I�8[�m�� �3f� �1x����������� *�<�N�`�r߄ߖߨ߀�����������WOR�`f�L���&�t� ������������ �(�:�L�^�p�����8������POd��� ��d���%7I[ m������ �!3EWi��DEV����� ���//'/9/K/ ]/o/�/�/�/�/�/�/��/�/?PALT ��81d�?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O&?GRI`f��AP?�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHo�OR�̀a �OZo�o�o�o�o�o &8J\n��������noPREG<>%��o�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~������$ARG_�L�D ?	����ӑ� � 	$�	+[�]�����ƐSBN_CON?FIG 
ӛ&��%� �CII_SAVE  ��E�<�ƐTCEL�LSETUP �Ӛ%  OME�_IO��%M�OV_H������R�EP�l���UTO�BACKt�0��FRA:\�c ���_�'`����=�� J� 	������ͿpĿֿ�6����	� 1�C�U�g�yϋ��� ����������ߜ�5� G�Y�k�}ߏߡ�,��� ���������C�U��g�y����a� � )�_�_\AT�BCKCTL.T�MP DATE.D;<��	��-�?���INI;0p�8�~�MESSAGT��^�_�ېi�ODE_AD��W�8�H���O�����PAUS��!��ӛ ((O ֒��
��*N< r`��������"����TSK�  ��=�C�	�UgPDT��\�d����XWZD_ENqB\�4��STA[��ӑ�őXIS&�U�NT 2ӕ`�� � 	 ����W�f I��M�b�����"9�(#>��T #M/� " Klޤ;�`� ��0}���c/�/_/�/�/�M[ET�`2�P�/�?�/<?�)SCRD�CFG 1C�`��\�\� 1?�?�?�?�?�?�?6��QX��??OQOcOuO �O�O O�O$O�O�O_�_)_;_�O�O���G�R����zS��NA���қ	�wV_�EDZ�1e9� �
 �%-��EDT-h_ʪ�_o�`/^���-��_��	������_�o  ���e2�oɫko �o�6k�o!hozo�o�c3Y�o��o�n���4F�j�c4 %��r���nN��� ����6��c5�a�>� ���n���̏ޏt���c6��-�
�Q��n�@Q�����@�Ο�c7�� ��֯��n���d�v�����c8U��_����0
 }~��0�B�ؿ�f��c9!ϑ�nϵ�  }Jϵ���Ϥ�2φaCR�oį9�K���߀�����n���zP�PN�O_DEL�_xRGE_UNUSE�_�vTIGALLOW� 1�Y~�(�*SYSTEM�* 3	$SERV_GR�R 69���7REGB�$d� <�9�NUMg��z��PMU�� 5L�AY�  <P�MPAL[��CY'C10����������ULSU��{������D�L�N�BO�XORIk�CUR�_;�z�PMCNmV��;�10��>��T4DLI�4�V���ߨ���'9K]oR�zPL�AL_OUT �Dcc�QWD_A�BOR��	��IT_R_RTN���Y�� NONS8�� �CE_RIA�_I��<FF_1�4e :[�_PARAMGPw 1�w�`_����Cp�  .� � �� � � � �� � � � �� � �  D�X $3!g-�<$��H$�T$� D*X � X "� B�kD1� 9X @� 6�?� <HE��ON�FIy���!G_Pv��1� �e �U??0?B?T?f?x?|�?�!KPAUSX�s1�UR ,Z� �?�?�?�?�?OOO TO>OxObO�O�O�O�OмO�O_�2O_�ey�PCOLLECT__�Y[ 4cGWEN��I�"cR Q�NDEOS�W���1234567890�W�S�p5b�_�Vy
 H�y)�_#oS��_oho T�AoSo�owo�o�o�o �o�o�o<+� Oas����� ���\�'�9�K����o��VQ�2W[ �� 9W�VIO �YcQyH&�8�J�l\��TR�2؍�(��
��j�� � ����%�_MOR҂!� + �'� 	 �5�#�Y�@G�}�k����Ӂ"��2?�!�!3 ҡ��Kڤ��$R_#�*_	�:Q:RC4  �AS yC  x�=A3!z  BC!�P�B/!�PC  @�*����:d��
�IPS$����T��FPROG %�*6߼�8���I����&RҴKEY_TBL  )V�R:P �	
��� !"#�$%&'()*+�,-./�W:;<=>?@ABC���GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~�������������������������������������������������������������������������������������������������������������������������������������������1��L�CKۼ3���STyA�д_AUT���O(��U�INDxtTD�FQR_T1_�Q�T2��7$����XC� 2����P�8
SONY �XC-56�9Q}����@���u�} ��А�HR5��cT0�B�7<T�f�Affrꬿ���� �������5� G�"�k�}�X��������������ǼTR�L��LETEG���T_SCREE�N �*k�csc:U$MM�ENU 1&�)  <��� y��Ã�= &sJ\��� ����'/�/]/ 4/F/l/�/|/�/�/�/ �/?�/�/ ?Y?0?B? �?f?x?�?�?�?�?O �?�?COO,OyOPObO �O�O�O�O�O�O�O-_ __<_u_L_^_�_�_ �_�_�_�_�_)o oo _o6oHo�olo~o�o�o �o�o�o�oI 2�X�hz���� _?MANUAL�ߕ��DB��L+�DB�G_ERRL��9'�� �\��n����NUML+IMK�d �p��DBPXWORK 1(�I�ޏ�����&�ŽDBTB_@ )��������qDB_A�WAY�_�GC;P  �=�װ�~��_AL��D�z��Y���M � �_)� 1�*����
�͏����6�@�_M&{�ISAЉ�@B�P��ONTIMJ�& ��p�ƙ
�ۓMOTNEND߿�ڔRECORD ;10}� �>�?�G�O����?��� 2�D�V�h���p���� ��*�߿�Ϛ���9� ��]�̿�ϓϥϷ�R� ��J���n�#�5�G�Y� ��}��ϡ�������� ��j���C��g�y� ������0���T�	� �-�?���c���\��� ��������P����� ;��_q����� (�L%�4 [�����^ t�l!/�E/W/i/ {//�//�/2/�/�/�??�/z�TOLEoRENC��B�ВL���CSS�_CNSTCY ;116�  ?Β�?�?�?�?�?�?�? OO&O8OJO`OnO�O��O�O�O�O�Oc4DEVICE 126� b�*_?_Q_c_ u_�_�_�_�_�_�_?��d3HNDGD �36�Cz�^LS 24]�__oqo��o�o�o�o�o�_e2PARAM 5��B��t�dc4SLA�VE 66�e_?CFG 7��gdMC:\e0�L%04d.CS�V�o��c|�r�"AM �sCH�p&a&�P�n��w��f�r�����ÀJP��>��\_CRC_�OUT 8U�����oEpSGN �9U�Ƣ��\��15-OCT-�22 18:03��p�02��4�:41�p9V UBu1�݁�nހ���o��Im���P�uG��@uV�ERSION ���V3.5�.11E�EFLO�GIC 1:ݫ 	6��|�C����^�PROG_E�NB����͢��UL�S{� ��^�_A�CCLIM|���Xs��WRSTJN[���ţ�^��MO��¡Zr,�INIT ;ݪs5᡻ *�OPT$p �?	i�B�
 	�R575�c��7�4��6��7��50��R�Ƣ2��6��X�>y�TO  ���t?�Y�VP�DEX��d���@W�PAT�H A��A\�E�����7;IAG_�GRP 2@�k�,�"	 E��  F?h F�x E?`�D���û��V1"�ü��XT0K�9�Cf�py�p�Y�dC�pqߪB�i�ù�mp4m5 78�90123456���;����  �A�ffA�=q�AةpхAʯ�HAĩp����~���A��Mk,���@��tp�p���W0A�T0T0�pBA4ü Qô���
����(�A�A��
=A�L����A��
A�Q��A��������e�����e� Pe��:��{A�d������dѩp�������A�������́�r߄ߖߨߺ�@�E�G�A@�p:�R�A5d�/��)��#
P�d�l�������"�4�F�@�Pz�A�J��c�?��9p��A3\)A,��A&����0���Ю�����@�cP�]�W�AW�P�J��UC��<d�4�-d�%G��(�:�L�^� @���$HZ�� .|����bt � 2Vh�x m�����[���s������=�
==�G=��>�Ĝ���7���8��b��7�7�%�@wʏ\"&�p�.%���@�Ah�p9 A���<i��<x�n;=R�=s���=x<�=�{~Z�;��%�<'�'�~ �?�+ƨC�  <w(�U� 4"w����&����%ùf��@?Œ?� ?@?R?g��$^?�?"?��?�?�?�?�?�?)�7L?S�FB$��/"Eͽ�>OG�ΐԬq��sD�5L4�x�CA��Gb�@tφ���-_7_�C���_;�/_�NED � E�  Eh� D[PbRD_¿�_��8�?�p3���}��C ����|�Q4|3��2�C,�{����QE P C��/GC�7�<�{_�_w_o�K:o@bù��Y7a,�5����6���?��o�o	o�o�o�o�o��oÿհCT_CO�NFIG ���Yt؃e�g��ԱSTBF_TTS�
ęVs3����
�iv[�MAU����Y�MSW_C�F*pB�s�!�OCoVIEW}pC�}���6�
��.�@� R�d�w�������ȏ ڏ�{��"�4�F�X� j���������ğ֟� �����0�B�T�f�x� �������ү����� �,�>�P�b�t���� ����ο��ϓ�(��:�L�^�pς��|RC�sDJ�r!ϐκ� ������7�&�[�ot�SBL_FAUL�T E���xu�G�PMSK_w��pTDIAG F.y��q�IUD1�: 678901�2345��;x�MP �o!�3�E�W�i�{�� �������������/�A��( W!�J�"�
��vTREC	P����
�����M� (:L^p� ������ �$6]�o�l��UM�P_OPTION_p�ގTR�r`s�ٝ�PME^u�Y�_TEMP  _È�3B�P s�A�P�UNI�p�au!�vYN_BR�K G�y��EMGDI_STA%��1!�rL NCS#1H�{ �K��9�/_}dd�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO��O�O�O�O�I �!�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXo�J O�o�o�o�o�O�o�o +=Oas� �������� '�9�K�]�wo������ ���oۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� o�]�������ɏ��� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�g�y��ϕ� ��]�ӯ������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� _�q�{�������� ������/�A�S�e� w��������������� +=Oi�s� ������� '9K]o��� �����/#/5/ G/ak/}/�/�/��/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OY/KOuO �O�O�/�/�O�O�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oQOcOmoo�o�o�O �o�o�o�o!3E Wi{����� ����/��o[oe� w������o��я��� ��+�=�O�a�s��� ������͟ߟ��� '�9�S�]�o������� ��ɯۯ����#�5� G�Y�k�}�������ſ ׿�����1�K�9� g�yϋϥ��������� ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�C�U�_�q��9� �Ϲ���������%� 7�I�[�m�������� ��������!;�M� Wi{����� ��/ASe w������� //+/EO/a/s/�/ ��/�/�/�/�/?? '?9?K?]?o?�?�?�? �?�?�?�?�?O#O=/ GOYOkO}O�/�O�O�O �O�O�O__1_C_U_ g_y_�_�_�_�_�_�_ �_	oo5O'oQocouo �O�O�o�o�o�o�o );M_q�� �������-o ?oI�[�m���o���� Ǐُ����!�3�E� W�i�{�������ß՟ ������7�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿��� /�9�K�]�oω��ϥ� �����������#�5� G�Y�k�}ߏߡ߳��� �������'��C�U� g��w��������� ��	��-�?�Q�c�u� �������������� �1�;M_�� �����% 7I[m��� ����)3/E/ W/i/��/�/�/�/�/ �/�/??/?A?S?e? w?�?�?�?�?�?�?�? O!/+O=OOOaO{/�O �O�O�O�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_�_O#o5o GoYosOeo�o�o�o�o �o�o�o1CU gy������ �o�-�?�Q�ko}o ��������Ϗ��� �)�;�M�_�q����� ����˟ݟ�	��%� 7�I�[�u�������� ǯٯ����!�3�E� W�i�{�������ÿտ �a���/�A�S�m� wωϛϭϿ������� ��+�=�O�a�s߅� �ߩ߻��������� '�9�K�e�o���� �����������#�5� G�Y�k�}��������� �������1C]� Sy������ �	-?Qcu��������� ��$ENETMO�DE 1I^�   � (/:+
 R�ROR_PROG %*%}/�)�X%TABLE  +h�/�/�/�'�X"SEV_NUM� &"  ��!!0X!_AUT�O_ENB  �D%#U$_NO21 �J+9!2 W *�u0�u0�u0	�u0(0+t0�?�?�?N4HIS3
 G;_ALM 1K+� �u< +�?/OAOSOeOwO�Or�?_2T0  +�s1:"�J
 TCP_VER !*�!u/�O$EXTL�OG_REQ�69�E9 SSIZ)_T�STKFYc5�~RTOL  
{Dz�2�A T_BWD�@�P<6�Q�8W_DI�Q L^G48$
?"�VSTEP�_�_
 �P�OP_DOh_!F�DR_GRP 19M)B1d 	�Ofo�: W`�������glpw��qŗ�?�I ����fWc��o�m�dAҔA�׼h�b���A�`Cm�o�`�c��A���bu�A\���o#�o �YD}h��@���A8��>��Β� 
 E㻀�c�p�r��C �B��8�#�\�G��C`}dC��N���B�{��F�@7UUT��UTF�Ϗ�j��s���E�OHc�EP]��O���#M��*�KA�����?�F��:6:N�r��9-�z�������� �YJ D�R�c ���|Z�����+FEATURE N^��P>!Ha�ndlingTo�ol � mpB�oEngli�sh Dicti�onary�
�PR4D S�tڐard�  �ox, An�alog I/O~�  ct\b+��gle Shif�t�  !*�ut�o Softwa�re Update  fd -c��matic Ba�ckup�IF �O��ground Editސ��g R6C_amera3�F7��Part��nrR�ndIm���ps�hi��ommon� calib U䗠�n����Mon�itor�Cal�M�tr�Rel�iabL��RIN�TData ?Acquis�Z��ϠC�iagnos���0�<�almC�o�cument Viewe�\���C��ual Chec�k Safety���  - B�En�hanced U�s��Fr���8 �R5�xt. D�IO �fin� �(�@ϲend��E�rr�Lm� D �p^���s	�EN��r.�հ �P�r�dsFCTN_ Menu��v8����m�FTP I�n'�facN�=�G���p Mask �Exc��gǱis�p��HT^�Pro�xy Sv��  �VLOAאigh�-Spe��Ski^ݤ ef.>�Hf�~ٰmmunic���ons�
!
���urE�'�7�rt� F4�a�connect 2;��Incr`�str�u���� Sp�KAREL Cmod. L��ua���OAD*�=�Runw-TiưEnv�� �D;�(�el +���s��S/W�.�{�Licen�se����
����o�gBook(Sy�stem)蔭�J�MACROs�,��/Offse�S�Z�MHٰp��� wj73ΰMMR���l�35.f��e�chStop��t��R� ize*�M�i��O� 2�7�xp��0����miz���odM�witch�����a�.�� v����Optm��4q9���fil���ORD��0�g�� �8496�ulti�-T������C�PCM fun�,��.sv�o�O���� �^�5�R�egi��r��	�!�2�ri��F�  �H59k�1�Num� Sel*�  7�4 H��İ Ad�ju���adiṇ�O� ,[���tatub��\У��������RDM Ro�bot��scov�e� �d emt(�ٱn� SW��>Servoٰs��ꒄ�SNPX �b��1��g P�L�ibr���1��ڐ 9� ɰ.�30g o��tE�s�sag� f�E�@ e����"g��/I_�
�I�TMILIB���� ?P Firmn��8�^�F�Acc����<0���TPTX����510.� eln����������H5�73�rquM�i�mula��� 2n�Touz�Paxъ�1� T��6���&��ev.��I?USB po�����iP�a�� 0\�sy nexce�pt��3 <� \h�51 ����oduV#��9��Q��VN�k"6PCVL�{&�^}$SP C�SUI�d���+X�C��auҠWeb' Pl���t? �# S��\"	2��������S�&ު�V?8Gr{idplay��`&� ��8�-iRb"�.� @ � R-2�000iC/16�5¦ d+�+�la�rm Cause�/1 ed�<0:�A�scii����Lo�ad��V4�3Upl8�0�_CycL�c��m�ori����FR�A[�am�) td=t��NRTLi�3�Onݐe Hel�ݨ 542*�PC�`ρ�4�`�]�1t�rߵ48��ROS/ Ethv�t[��n�10\ҠiR}$�2D PkߵDEaR>1�E����of�AX��ΰ�FIm��F���� z��64MB DRAMު�@:�9R�FROA[�Celal3� ����shrQ�
��Zc���ÍUk�p�� pide�WteyL�s��|0\z��!CtdѰ�.��@"E7mai��li���B+�\�� R0�qZ$�GigE�N�4OL�@Sup"��b�W38oa�~�cro���� ��4��QM��Fauest�A>�j�� �miH9.dVirt`��W��0{&ImM��+T���}$Ko�l �Bui��n�յ'A�PL�&��MyV6� �"�0�*CGP�l����{RG�'p�{SKBUW�RQ�)K�&cm\:��z��fX�)�O�võ(TA�&spoҠ-�B�&��
 �I�\E P�+�CB�'fg-��&"k  �E��sv�b���vv�3��S_k��TlO;-�EH�f6.
��E�vfx_z�)�V��tr>�)�hZ%.�F�& � ��r���*�G�&���њr�����H��РJzCTIA2c�pw4�LN�1�Mr�" #[��g�""�M�-�P2�~�T�@����vxui$�-�S�&�S�&�*z4�W��2.pc�)wVGF��fxwʪ�VP2AU \fx���N�if�u���w"in��VPB����)��s�D��*��a<s�F�5 M״�s�I��c;�{&Traİ���U,p  ��<���2��RDp	�N���HY���p��-���H���Øp)����� �ϭ�����ħ���rд�<���í4+����'9L���ӎ���y�9ӫ�c<3�U��B�O�q��u��kߍӍS�y*�ߩ�\Yy<����k�W����τ�Yx����:��	������<�5�o�e/�Q�ψ�,�K�m���g��^~����u�2��A���������F��<����y�)����|����1�m�.y�+�M��8G��i�7n��c���1籖 ����yW�����7�{�����6�Z�������uk��[�|��!��?�ϔ��9iB\����_�#�{�x@.��wrst���B�� H68��@�H)T@J�EENsDI?��tql[}
_�w�P��TQ (��I)# "���PA���8T�/��85/A#bs;/�C/U/�,q �/B�Gp�/�#��/�"�36�5�R ?!2e'pai?5!:/Y48W���%INTo?e?�_.q�?4)��?�2p�a2g�?�F O��?A�ad6?��t <ZUD2gunOOqCG533R?�D�0u�O�/�Mcm���OO�LNT�?��P_�Ĕ�`0_QR7�L_�Cfi._pH?_,_f'R50�_�SAF-F�_�7�w.vo��_�_8�/�dM Cbo��̜o�bvrEo��pa�a�oaD�@�osF-AS-sS�p'Isq(�PCesXPL�O�tlo_�ut\a��Oh%afvh%- B��/����C�$��srp�?@_�?`Dw�}�bA�����h�`௏]T�ˏ�sgc�h�os�t��CG\�s;��us�?���S9g�/�G J�����GDǟi$"�o�g3diʏ!�fd����?h%J64S��Tut�o�O�?s����F�_ ����E�0���D`!�)�NO4E�O�i$3II���iwjOl�`ž��>�?*�lb
��V��vjr/��
����7��ϥ�_�?zG7\2O�EG��Ϲ?���01� ޯ��_d�oi�A8��c�50�>�x����"Lo�h%����dj9�﴿ƿؿ��c� up9�C� j�9{�E��L��Ek,B串����oS_e_��&/��O}�j94JϬ�duZ��U���=d;�����8���r7�Dhu���;]m T��������2f�a���M�`���P�-4r V���O" #S�dw�c�P�in�`�ḁ?& HTuReLf���
�?hc��g�r"��q.JG"�erM/��/ �/�LRA^��uH71��/�tCK�/<eTX�P/?i�k1/m5k.�f��riR�eH1G�/�/ cr�NNHGRf?L�iY�d7�hOuX��H\mO ��oρ�;H��DD@�O ��*�<�:I�?�?��dϜR�_ hd�gh�gOO�_���gmh�_h�m��XO�o|O�O �o�O\/�o0�f�gm�o`��`e۠;iov��yt��"��u�R60���#tm�o_�#1��fdr,op7��_����lp>oh���O�~ ߏ�d&gts���&dޏ�/`�o�o
�J?<�vrF����v.R���Ɵpld�56�%4�0/����reeK�m�XP�)�KCO*O|%56 ?�OZ� o~����E$�io����jߠ���l� ����OR��LO1Fvod��_IF��$� � ߪ�DߦX!B� U3ce��t�4 ���(M�O�5)e?Ƕ/����1?Q�D�uk �'�|����`�boto�����-���6�p�0eS ��on*��� ^�lB'����Տ_�q��_�rdk��4f�� C(ҿȿ¯ԯ�������̟�����
I���571��t�a3di39Tar��lփofk�������vP�a�@� PJ��|*��������3et�4epg���e�d�� E�5�R�I  Hw552� 747��21�pWel�R78�,� �0�ETXJ61�4��ATUP�  wmfh 5#45�p�"6�pk��VCAM  �7\awCR�I@ ED" G U�IF)!28  =j�CNREM�`��63�a�SC�H  4C D�OCV� CSU�i�!0 D s�EIOCE�54��#R694 we!!ESET=S#!3!��a 73!fanu�MASK���PRXY�_"78� �0�OCO��"�3=P[�#"�ER �J�" 7�!!J7�74#!39�  Eqq�G1�LCH 0�#OPLG%J5y000#MHCR)%sPS�17#MCS �4D"�04 O#J55< [#MDSWe!Y13MD#1s#OP#1#MPR$07�0w"0p�#�  �#PCMX �#R0A�#� &�0�0�#� ( �&0�$590( �#PRS� 3�J6903FRDz@ 02RMCNy�7ndM�93 �SNBAA�8�00�@HLB  �"Lo�SM�A0� (Ww"4 oni�t#!2  II)��TC [#TMI�Le �B�`0"K3��@TPA� �QT�Xa�t\j�@ELL�BM250`0/D8�v�$78�mon�1�95d SD95\FU�EC 0OP� UFR(@ ��;!C@ \�@;!uO�0pt"VIP�@�#� I�@0�!CS9X� �#WEB �#wHTT \stB�24 �#CG�Q#I�G�Qtopm�PP3GS!��PRC�@S#H7���w!6( �8��![�R RBB-� Ci�B01rog�w!#IF#"098`-!!` �@�A64�(AaNVD�!Ld�1h 6a68( c�`d �SR7c!te.p� 0kaч@�bc`� �CLI$0?�sb$c9�G MS�"5a�` -� A� STY�@a;l �@CTO �CwJNN0J98��ORS�0G��b�g� J�`OL�1Ab�n: SENDu�to�!L�Q���@*r#�SLM� 8�"FV�R� MCHN0CSW!SPBVP�� KPL� ds �qV$0��cCCG $p�aC�R�0
Np�QB� 8�7.f�QK� j7a0*`�p�0'3CSq7Too�CTQ��&�qTB�P�N��@In;pqC�@�Q#�� �p,#�p ��. %��$07#%� `8D#TC6� QSQ"TE� [#Xm� �tTE� gt"m�P�TTF�Q[����@�#CTG�Q�"����@�#CTH `�TT�I�@#CT'Qeqs�PCTM�@SC��$0gS��0bodyzqP�@  ���� �1� d��q�aus�a9��P�[�qW `@06; GqF `8�V@VP2@ G623R i��@j?��g� `n�g�B `"D g�D `��g�FX wmna"PVPI���+ G V�!#V	` 7 23�RVK�@Np��@CV�Q31�9�34.�vo R�erne땗��$��i��r��땁h���A���3�7� ��"�\srv����b�3b�/- Sr�B"0��<�A�J935땿B^�5 (S�O�� �g �1�1�R�|�j93땷b��E�N�5�� awm��SK� Lib �������� ����	 �"|�h��h�#��b�wmsEk�nE����q�6��pyE�  ����!�02�t Fu�ïբ6ۯm��ujKi-�I&���8k� �8!�Ń�땼P��2�2�2�Mai'�on��_�/r�;pڦh;�;�G��_r���!��4\ֶORCt��+�5�� "T¦aTP��hQ�652�a1��4���<�xk��(���ߦ�t�P��Q�rֶSB�� ch_ ����)�t!0�B�"̿ h�h땇�;���c� �����������>�<�Rp� \toֶ3�F��cl�W��2p� "���������� F����b� Qt�a�ϒ�0t��ܐFsȒ�7�6�p�t	� Ad���582��ob��|*{�\a���FMQ ���A�mcigֶ�I�or�pwI�j�rfm���Fc���@1�EYME~� w���R��b�4�K2Х70.�9E�ld,�C�6� 1PTP]��\�.�"AD.�F�p&3 k���ask�D�ȍ`4���۳dֶ�ے��ER~�7 R �ƫ/�T�?)�e�rv�G?Y?k?}?�?�?ӹapa��	d�Ъ��r�4�M��teD����79!J�d/�2��G�p�ac�T� �<6�b�/� QO��$vc>�,@Vg�����eYW��5/� 1BJ�h���R5:�d���0�@��I_��raj��e��he(}�$`��5(Xa�@���et榻�1Otdj���,�_h�\	UI�/k�jo�FO��`^�°�F��r��qW65�q���K �'6ڦus W'�b,'��'?:��n��MFR��;�]�lf�ǯ�fr>֛�w�p�/�,� �_U[ǀ�мn�x'_ i�{�����O���pJ����[@�o�in7L��O�9�\^� � R����+m�i2״h �j��҇-� f�nt >�M�A H�I  �H5529� �(Cߑ21��leR78�c�ߒ�0AcaJ6�14���0AT�UP�����545.�t-fl�6yE=��VCAM�tFLXCRId���o�wUIFULX ��28��mo�NRE�u'��63��WQ��S�CH��Cn�DOC�V�gϠCSU1�c�xr�0$�;�EIOC%tx\cF��54�oQ��9T��;�ESET�Tem!o?�S�/��7S�{�oMASK��70���PRXY�T�`��7t��`�OߐOCOe��\?�3�ô`>��0�{�?��|�-��o7n G?�39!'ߑ�õ H82L�CHd��@IOwPLG�tCGM?��0��GЎ�MHCR��Go�S�/1_�CSn4�cgm��50T�ě?�5$�[���MDSWMf.�D�����{OP��X/2L_�PR��K�����{��n�883n�CM��/0iA,��0�Ő`z~�5#�\h88� ��+�?�D���.?����4��0D�3��o�S�4����9��,i�FRDd�/2E�/��MCN5�H9y3�K�SNBA�U�"R��HLB��S�M�՛ñ�T���J512�SaߐTC4�\�TTMILe���P���A|�TPA����TPTX��5N��TEL�ԫ�0��P��8�˳���K��95����95��8�88��UECd�r;t �UFRd�_�_�Cd�2e-�VC9O4��VIP�;���I�TAX~�CSqX�����WEB4����HTT4�ka���2T�2M/So�G<#��QIG��< �.�IPGS=t\r�xO�RC��aߐ7��/a��6D�s@>�R7#��!��Oq�Ҥ� �P��Ҷ;�A���KÑ�.$�0 "��4�����NVD4���#�Ad�ap��8D���68�����R7���P��D0��a��o�bܠ. 7CLI��l\-C���CMS�'��4�wd "ްSTY�n[�CTOT�tl��sNN����ORS4ĸ;�1 ��ltiΰO	LS�( E���0�TЊ��L��6�@���9�@ ��LM4�HV� o�VR���CSshc>�PBV�4䫁/�PL�
AP�V��ust>�CC�G4��0nCR�4 H5��B���=K�H573���x?����\cms�n#�st.~TB��P�! ��7�C��x��?"�awsh?"���I0?"��3�T�Cd�K�A 4�\sl�"EĤpP��� 4�C[П"Ԥ8c��"4�(�.�CTF��c��"����CTG�73�m#G�THd�hd� �I��K�CTC�;59m�CTM�5�M����Q0��re\g�P���12�@�04�����%S��13MCTWd�9l[@_�GFd�SE]�P2d�t+��2�ա ��2d�ell��PBd�I���1Dd��a�1�F��tap VP�Id���CV�!Vtq��UA��CVK��ۣCV#�coreAL���H"�Hp!8�HK"�Hatc�J$�H�4�I� �IL0H�I�2�H��H+2�I�L�Y4=�H���Iec\a�I�2 Z93�I@{�H�@NZ+��H 1�F�K48�Z<A�Ht{@�Il �Z;"�O�Fs\! �Hk"�H{"@o�F[�PZ!o�Z���J��Tok���H��H\��Il�Z���Z2=[ng-[gToo�I�p�j(�nj�robt_�Xbt1.�JL� iur�o�I@��i�!��F��POz�ling�j��y���Y"r^zۢ�I�p��Geat^j�]��Z��_je�����_��lkҠHm,��H|��Zz��A�I  �_��  ���Gvhm��J{�svnj���H4�9\�J�@L�Ij7�49{P�Zt\j0Nj�@_"g.pjmgcal�0�fu�J��^zhm-��_bg����o�\ͫ �1�H!� j��;����MT "�(Cu�zk��&bgft�JlpX����GCT"���Gfc<]�˝26\fߟ�926�l\� Ίu��>m��;�Mul?�Q��7\^�K����7-[˝���_�61nNj48.� H- ԠH�@R_�L^ziPae��K�Я�F8\}��}�����Ћ� � R<k,�ticMoj+@�OoQxs-@�"�3�C�S j+}LB-[5s HNj+� co~��L��z��f�k˝lb�jll����-˜��k/�.���LЎ�ki;pJ/�on,�J\A���8�SK"�� ��uto�o B�������kwm� �o��Htp�ʜ n}F��ex-�˝��x��J�a^jlL�je����i��a��/����rej�1X�o�Vor�zR�ߎ��e T�Z[��[l#clN��߭�SOžgGZD��to�{�+B�H643N�`�S1G/o��sg�a�Utui��;`�J���`�;�ndm�ndiN�{/�/�/�/�/�/ �/�/??/?A?�?���riΪ! -Kj9�50/�n �zk]8c95n/�O�t �Z��wsg�K,�>��wiag� SGJ�Ю�ogu���KO�]Ltw>_@	J64t�1�s�{F O>�F�cdݛ��`3_���r-��N74�y�-�3��RINnzlly��(m^���L����sgc�zI" �#?
+�oߡ\tw /��0.�@�"���f��_�[y�Kmm�K}d�ct^�t]�+�
P�RZWCHK
kA,�;;`y<p��lK�t��LN*R85j� �@_jR ���t�iN�g WJhe�cN�L�F����wl�Z|*�dat��ʛ�greN��o�  ST�D�r7LA[NG�Aoc�e�`���Q�7��R8�70�{��8 (=P�ogge���!�58\�P�ATTs�� �t\���c "B�@Vx��1�patd���O���������{q㕔�5�a�p[�m��\㕻�7�\aw ��@�a��p6���x��ϯ�gmon���d��0�B�m�;A���\ ö��K�I�M�HCR�51 H�����g\o��@��R]� H54ۿm�<@�E���;!�����o#mm�;a��R�|�N㕬0F�C��W�P�)Ai6�� Fƫ�{�.�itx�#{ ���iaio����De�6�eve����72� R�@RƜPg��a�dl��nt��K�RBT�tOwPTN`772'�CTK"'�g�(䔠<�)� "AZ'�;q8'�q'�tzn&�{ �E'�Ama��- �Mu��ncInDPN����Ҟ��872��|�d��(��������#����masy��y �"M��o��䃲��et����\p1�����d\ ��f���lZ����lp���9���`��8+ V��ail��?� �䇢�䓢��zd�<��k`��73.f��iwrdg��- i���e\ ����� S0.j�021"�1W ��p(�`�4�� (i��e,"� "���+�^��core_�I���l`F��AY��AB���@����H�����AwBIC��Par;�M�ai������<�v c\�ITX>����  ����1���g Jcl;ib��ShiW�x4�� t994\��VSSF��� tt�\j9�f "O��w� t��$%ini�/��pٰ t�5G8�&,� t\vsR&x��L�%w� tamcl<S/+ref.�%#� tj��%m�� t[A΃&4\z�/�,z_�v�%A�%�a�%_o�l6��l% �%en	d�/<c?.?@?R5�o[?m>�6�/�dsh9f�/+trt�?<xOAE�'F  !�G0��$%��5vi�6���6 J92�F3��%O25 (�%�@e&�P�%k�4O dnw�zF��T�&`�XEpn��&g��? nw\nL�?�,nd�V��N;XfnF j���%se�V I/
&�q&фU���5r w�%/F�� �F�_�rclR&0X\pw/Y�90�Eo`t/"5Of "U//A+dprm�%g¨%��Xrsu/kmS�T_ L`�6/OŔpM�LO�j���nO1|h�ODnopn�|YCwrpR/��l���E<�Pe\ga<��Krgas�o�k���f�v��4xt�f�?m$ra�o�la`0�omk�_�TamN6�+�4�`'9K0.v �Wې�%�@�Ft��XE� sV��ДJ73=7�%|*�%,P̲�hB "+��Kwc�fF& I����99�8�vtomzFut vV�_	o;�YC��F�:8\F&�Y/� 0:��f��deb^V���$�0zFؠ"��gL���<9\�&��9�W�r}  �su"�st��G��X �f� U (�fagn�F PzFϜ6�Via�TX����vd��w��g��HzF7- O�W CH� ��$723�F���E( A�ÿտ2蚽Wc��W�svF& S�W�JRi6��_�RVo RV0���ӊ��vt�MG\etF�XoN�o�FAr��x���+�1T�F�?teR� J58��O  34	Wgl�e,�%,�j�Dq\t0"��zFwIta1lU#TA�VϜ�gw韗M�ad�W�Oa���6d� M��e�FT��9�0 H�%NT��R�69������ir�\ʆMIR��ӊenʆv���F|�3��I'TCP��Ta0�p���(MM7G�eT�o/ \tpʆI��YB'busJ׈�m��I�@zFȀ��F�����t/��W�'g, ��4`R_(!sw�&s_YC�67\JF��Tf_����Dfw��W��4gachg��a96_�d�� _���_rV��% 99�YA�e��$F�EAT_ADD �?	����~�  	�$ YA//%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /�A�S�e�w߉ߛ߭��������DEMO� N�   ��*� �2�_�V� h������������ ��%��.�[�R�d��� ��������������! *WN`��� �����& SJ\����� ���//"/O/F/ X/�/|/�/�/�/�/�/ �/???K?B?T?�? x?�?�?�?�?�?�?O OOGO>OPO}OtO�O �O�O�O�O�O___ C_:_L_y_p_�_�_�_ �_�_�_	o oo?o6o Houolo~o�o�o�o�o �o�o;2Dq hz������ �
�7�.�@�m�d�v� ������ƏЏ���� 3�*�<�i�`�r����� ��̟����/�&� 8�e�\�n��������� ȯ�����+�"�4�a� X�j���������Ŀ� ���'��0�]�T�f� �ϊϜ϶��������� #��,�Y�P�bߏ߆� �߲߼��������� (�U�L�^����� ����������$�Q� H�Z���~��������� ���� MDV �z������ 
I@Rv ������// /E/</N/{/r/�/�/ �/�/�/�/???A? 8?J?w?n?�?�?�?�? �?�?O�?O=O4OFO sOjO|O�O�O�O�O�O _�O_9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l���������Ə ����)� �2�_�V� h����������� ��%��.�[�R�d�~� ������������!� �*�W�N�`�z����� �����޿���&� S�J�\�vπϭϤ϶� ��������"�O�F� X�r�|ߩߠ߲����� �����K�B�T�n� x����������� ��G�>�P�j�t��� ���������� C:Lfp��� ���	 ?6 Hbl����� �/�/;/2/D/^/ h/�/�/�/�/�/�/? �/
?7?.?@?Z?d?�? �?�?�?�?�?�?�?O 3O*O<OVO`O�O�O�O �O�O�O�O�O_/_&_ 8_R_\_�_�_�_�_�_ �_�_�_�_+o"o4oNo Xo�o|o�o�o�o�o�o �o�o'0JT� x������� #��,�F�P�}�t��� ������������ (�B�L�y�p������� ���ܟ���$�>� H�u�l�~�������� د��� �:�D�q� h�z�������ݿԿ� �
��6�@�m�d�v� �ϚϬ��������� �2�<�i�`�rߟߖ� �����������.� 8�e�\�n������ ��������*�4�a� X�j������������� ��&0]Tf �������� ",YPb�� ������// (/U/L/^/�/�/�/�/ �/�/�/�/ ??$?Q? H?Z?�?~?�?�?�?�? �?�?�?O OMODOVO �OzO�O�O�O�O�O�O �O__I_@_R__v_��_�_�_�_�_�_m  h$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ� ����0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲�������|���  � �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p�� ����� ��$� 6�H�Z�l�~������� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ����������	�,�>�P�b� t����������� ��(�:�L�^�p��� ������������  $6HZl~�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o�i�$FEAT_�DEMOIN  �d�D`�`�,dINDEX9k�Ha�,`ILECO�MP O���zaGb'ep`�SETUP2 �Pze�b� � N �amc_AP2BCK 1Qzi?  �)h�o"�k%�o`}` Ae�om�o� � �V�z�!��E� �i�{�
���.�ÏՏ d��������*�S�� w������<�џ`��� ���+���O�a�🅯 ���8���߯n���� '�9�ȯ]�쯁���"� ��F�ۿ�|�Ϡ�5� ĿB�k�����ϳ��� T���x��߮�C��� g�y�ߝ�,���P��� �߆���?�Q���u� ���:���^���� ��)���M���Z���� ��6�����l���% 7��[��� ��D�h��i�`P��o 2�`*.cVR`� *c������JPC���� FR6:D�.�4/�TX` X/j/�U/�,;`%/�/�*.FM�/�	��/<�/<?�+STMG?q?��]?"�=+?�?�+H�?�?��7�?�?�?EO�*GIFOOyO�5eO"O4O�O�*JPG�O�O�5�O0�O�OM_�JSW_�_�� Sn_+_%
J�avaScript�_�OCS�_o�6��_�_ %Cas�cading S�tyle She�ets0o� 
AR�GNAME.DT_o��0\so1o�Q�d�o`o�`DISP*�o�o�0�o7�e�)q8�o
TPEI?NS.XMLg�:\{9�aCus�tom Tool�bar��iPAS�SWORD.��FRS:\�� �%Passwo�rd Config@���������� �r�����=�̏a� s����&���J�\�� ������K�ڟo��� ����4�ɯX������ #���G�֯�}���� 0���׿f������1� ��U��yϋ�ϯ�>� ��b�t�	ߘ�-߼�&� c��χ�߽߫�L��� p����;���_���  ��$��H����~� ���7�I���m���� ��2���V���z���! ��E��>{
�. ��d��/� S�w�<� `�/�+/�O/a/ ��//�/�/J/�/n/ ?�/�/9?�/]?�/V? �?"?�?F?�?�?|?O �?5OGO�?kO�?�OO 0O�OTO�OxO�O_�O C_�Og_y__�_,_�_ �_b_�_�_o�_�_Qo �_uoono�o:o�o^o �o�o)�oM_�o ��6H�l� ��7��[�����  ���D�ُ�z���� 3�ԏi�������� ßR��v�����A� Пe�w����*���N��`���֦�$FIL�E_DGBCK �1Q������ ( ��)
SUMMA�RY.DG�����MD:3�s����Diag Sum�maryt���
C?ONSLOGi�L��^�������Con�sole log�����	TPACC�N�R�%:�wς��TP Accou�ntinρ�F�R6:IPKDM�P.ZIP�ϯ�
����σ���Exception ߱�_��MEMCHECK�m�Կb����Me�mory Dat�a��֦LN�)n�RIPE�\�n����%�� Packet L�κ��$SA���ST�AT�����ߋ� �%�Stat�us��<�	FTP�����r�����m�ment TBD���� =�)E?THERNEU����B�S�����Eth�ern(��fig�ura߇���DCSVRF���������� veri?fy all٣�M(��DIF�F����/d�iff�PB���CHGD1�x�� �FQ&���	2�� q5�YGD3�8��'/ �N/��UPDATE�S.m S/��FR�S:\k/�-��U�pdates L�ist�/��PSRBWLD.CM�/«��"�/�/�PS�_ROBOWEL<1���:GIG�ߊ?�/�?��GigE� ��nostic�*�ܢN�>�)>�1HADOW�?�?��?5O��Shad�ow Changye��٤,8+�2NOTI��O"O�O���Notifi�c��\O٥O�A ��_��2_կ?_h_�� �__�_�_Q_�_u_
o o�_@o�_dovoo�o )o�oMo�o�o�o�o <N�or��7 �[���&��J� �W������3�ȏڏ i�����"�4�ÏX�� |������A�֟e�� ���0���T�f����� �����O��s��� ��>�ͯb��o���'� ��K��򿁿ϥ�:� L�ۿp����Ϧ�5��� Y���}���$߳�H��� l�~�ߢ�1�����g� �ߋ� �2���V���z� 	���?���c���
� ��.���R�d�����������$FILE�_� PR� �����������MDONLY� 1Q���� �
 �)�@_V�DAEXTP.Z�ZZ��p�G�L6�%NO Back file !��U3�M��7 ����G�&�J \����E� i�/�4/�X/� e/�//�/A/�/�/w/ ?�/0?B?�/f?�/�? �?+?�?O?�?s?�?O �?>O�?bOtOO�O'O �O�O]O�O�O_(_��?VISBCK����>*.VD)_s_��@FR:\BPI�ON\DATA\�^_R�@Vis?ion VDt�_ �O�_�__o_Ao�_ Rowoo�o*o�o�o`o �o�o�o�oO�os �@�8�\�� �'��K�]����� ��4�F�ۏj����̏ 5�ďY��j������ B�ן�x����1����ҟg���MR2_G�RP 1R���C4  B�O��	 
������E��� ֯�r���O�HcEP]��O��#M��
�/KA���?�&��r���:6:N{�R�9-�Z���A�  v���B�H��C`}dC�{�N��B�{���r���пὫ�@UUT��U����/����>��>c���>rа=ȫ��>i�=����>����:���:��:�/:6)�:��~ϗ�2ϔ��ϸ�������z�_CFG {S��T  ��a�s߅�0[NO ���
F0�� ���/\RM_CHK�TYP  ����O����������OM���_MIN��L�������X��S�SB7�T�� ��5�L�,�U�g����TP_DEF_�OW��L�����I�RCOM�Ѝ��$�GENOVRD_�DO��	��TH�R�� d��d��_�ENB�� ��R�AVC��U�UQ �Υm�X��|��q������ � �kOU��[��O�����⾥8��:���
,.  C�x �h�������B�ϡ�����\n�!�SMT'�\.����+�w�$HOS�TC7�1]K[[�Y� 	MM�MI�}�e���� /*��1/C/U/g/��/ 	�anonymou�s�/�/�/�/�/?  L^pM?�/� /�? �?�?�?/�?OO%O 7OZ?�/�/O�O�O�O �O? ?2?D?FO3_z? W_i_{_�_�_�?�_�_ �_�_o._dOvOSoeo wo�o�o�O�O_�oo N_+=Oa�_r �����o�8o� '�9�K�]��o�o�o�o �������#�5� |Y�k�}�����ď� ������1�x��� ��J��������ӯ� ��	���-�?�Q�c��� ��Ο����Ͽ��:� L�^�p�Mτ����ϕ� �Ϲ��������%� 7�Zϐ���ߑߣߵ� ��� �2�D�F�3�z� W�i�{��������� �����
�d�A�S�e��w����/ENT {1^�� P!�.��  ���� ��*��Nr5~ Y������ 8�\1�U� y�����4/� X//|/?/�/c/�/�/ �/�/�/?�/B??N? )?w?�?_?�?�?�?�? O�?,O�?ObO%O�O�IO�OmJQUIC�C0�O�O�O_�D1 _�O�OV_�D2W_3_�E_�_!ROUT�ER�_�_�_�_!�PCJOG�_�_�!192.16?8.0.10�O�C?CAMPRTGo#o�!7e1@`noUfR�T�_ro�o�o��NA�ME !��!�ROBO`o�oS_�CFG 1]��� �Au�to-start{ed��FTP��~q���F��� �����9�K�]�o� ���&���ɏۏ��� ��Wi{X����o� ����ğ֟������ 0�B�e��x������� ��ү�������Q�>� ��b�t�������q�ο ����9���L�^� pςϔϦ������� %��Y�6�H�Z�l�3� �ߢߴ�������}���  �2�D�V�h������ ���������
��.� @��d�v��������� Q�����*<�� ���������� ����8J\n ��%����� EWi{}O/��/ �/�/�/�/��/?? 0?B?e/�/x?�?�?�? �?�?/+/=/�?Q?>O �/bOtO�O�O�Oq?�O �O�O_'O(_�OL_^_�p_�_�_(�`_ER�R _z�_�VP�DUSIZ  j9P^S@��T>�U?WRD ?EuA��  guest3V$o6oHo�Zolo~o�dSCD_�GROUP 3`�E| Iq?YM ��nCON�nTAqS�nL��nAXP�n�_E�o9P�n�RT�TP_AUTH �1a�[ <!iPendan�g�~@}9PJ�!K?AREL:*���}KC����p�VISION �SET�`E��I�! \�J�t��s�����������Ώ��-���dtC�TRL b�]�~�9Q
@-F�FF9E39�D�FRS:DEFA�ULT��FA�NUC Web ?Server���� bvodL��'�9�K��]�o��TWR_�`F�IG c�e��R���QIDL_CPU_PC�9QB�@� BHǥMINҬ�a�?GNR_IO�Q�R�9P�XɠNPT_S_IM_DO�!��STAL_SCR�N� �y�+�TPMODNTOLY�!���RTY8��&�\9�hpENBY��c�ƣOLNK 1d�[�`�����1��C�U�ͲMASTE����&�OSLAVE e�_˴jq�O_CFGsϦ�U�OD��Ϩ�CYCL�E�Ϧļ�_ASG� 1f���Q
  W�9�K�]�o߁ߓߥ� �����������#�_ˎ�NUM�S�b�U
���IPCH��j�O�_RTRY_CN���Z��U�_UP)D�S���U ������g�θ`��`ɠ�P_MEMBER�S 2h��` $�e�>��Hyɠ�SDT_ISOL/C  ���r�\�J23_DS���q���OBPROCܶ�%�JOG�d1i��89Pd8��?�.���.�?�?�?OQNs��@V����3W~�����������PO�SRE��$�KANJI_m�K�i�p?MON j�k~�9Ry����//H�^�r��k����9%Th��p_L�I�l��kEYLOGGI�N���`����U��$LANGUA�GE ������ �!�QLG��l�q�9R��9Px�p�W  ��砬9P�'03X�k����MC:\RSCH�\00\��� N_DISP m���DAMK�SLOClw�آDz ��A�#�OGBOOK n���9P~��1�1�0X�9O%O7OIO�[OmN�Mɱ���I��	�5Ib�5�O�O�5��2_BUFF [1oؽ�O2A5 !_�2��=_?7Y_k_�_ �_�_�_�_�_o�_o :o1oCoUogo�o�o�o��oe4��DCS }q�= =��͏L �O-�1CUg���b�IO 1r� ��s20��� �����1�A�S� e�y���������я㏀��	��+�=�Q�|uE�TMl�d���� Ο�����(�:�L� ^�p���������ʯܯ�� ���7�SEVt��u={�TYPl����z�����!�PR�S���/S��FL 31s�}���π$�6�H�Z�l�~ϯ�T�P� l�i��=NG�NAM��A5�"e4UPSm0GI��\!��}��_LOAD���G %u:%P�LACi�2�3�MA?XUALRMI�c�8W�T���_PR�����3�R�Cp0t��9�M���3Eݗ���Pw 2u�� �1V�	i�00��� �߭�1��.�g�x U���������� ���8�J�-�n�Y��� u�����������" F1jM_�� �����	B %7xc���� ���/�/P/;/ t/_/�/�/�/�/�/�/ �/�/(??L?7?p?�? e?�?�?�?�?�? O�? $OOHOZO=O~OiO�O�K�D_LDXDI�SA����zsMEM�O_AP��E ?=��
 b��I �O_"_4_F_X_j_|_~R�ISC 1v�� ��O�_ ���_��_�Ooo@o�_C_MSTR w:�~_eSCD 1x�M�4o�o0o�o�o�o�o P;t_� �������� :�%�^�I���m���� ��܏Ǐ ��$��4� Z�E�~�i�����Ɵ�� �՟� ��D�/�h� S���w���¯���ѯ 
���.��R�=�O��� s�����п����߿� *��N�9�r�]ϖρ����PoMKCFG �ynm����LTAWRM_��z����и���6�>�s�M�ETPU�ӫІ��viND��ADCO�LXի�c�CMNT�y� l�g` {�nn��-�&�����l�P�OSCF����PgRPM����STw�{1|�[ 4@�P<#�
g��g�w� ��c��������� ����G�)�;�}�_��q�����������l�S�ING_CHK � |�$MODA�Q�}�σW��#D�EV 	�Z	�MC:WHSIZ�E�M�P�#TAS�K %�Z%$1�23456789� ��!TRIGW 1~�]l�U%�\�!�S
K.�S�Y�P�69"EM_INF 1�� `)�AT&FV0E�0X�)�E0�V1&A3&B1�&D2&S0&C�1S0=�)A#TZ�#/
$H'/O/�Cw/(A/�/b/�/�/�/? �&?� ��/�?3/�?�/�? �?�/�?�?"O4OOXO ??�OA?S?e?�O�? �?_CO0_�O�?f_!_ �_q_�_�_sO�_�O�O �O�O>o�Obo�_so�o K_�owo�o�o�o�_ �_L�_o#o��Yo ����o$��H� /�l�~�1��Ugy ���� �2�i�V�	��z�5�������ԟPN�ITOR��G ?�k   	EOXEC1���2�3�4�5�� �U7�8�9��� �������(���4��� @���L���X���d���Pp���|���2��2��U2��2��2��2ŨU2Ѩ2ݨ2�2���3��3��3(�#R�_GRP_SV �1�� (��>�>����O�b�"⸿�.�RƮ_Ds����PL�_NAME !����!De�fault Pe�rsonalit�y (from �FD) ��RR2��� 1�L6(�L?����	l d��nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲�����B2]���*�<�N�@`�r����<�� ��������,�>�P��b�t�����BJ�  �\  ��  ��  ���  A�  �B��T��� 
��������  �������B��p^���  CH Cѱ�P Ez  E��� E�` EE�;%��Z�*� �  �E��F�@V&��T Ai� dx�H�x��	$Hxd�d���}`(d� �8(xx$$�y Xtd D (DDdpWw X��	X�vXH�X���/y�y (� !��  f7%E	��Em��Xw$%XH$%P�� �/�/�/�/�/�/�??+?=?O?a?s=F�r?�?�?�?�6���E�#bE_�]��2  ذ���  ���?Kزd �3��(O:MO\OjG�0��|MTCҷ'4 � W%�O|�O�N  �H��O�JA  A��C�����_�OC_9W�
  � TB�LY��
��_�\�@Q�Y=�C�و�V�`HR0� ʒ_P( @7%?���a�Q?ذaر@��6�&س��2n;��	lb	  ����p�X��U�M`��X � � ��, �rb��K��l,K���K���2KI+�KG�0�K �U�L�2o�E	O�n��@6�@ t�@�X@I��b`�o��C�N����
���}v��#���` q�m�|�kQ?�
=ô��  �Hq�o`!b���9�  ��a� �B ���ذa�s�G��}2�m��o�q��v�O���E	'� �� 0�I� ��  � Q�J:��ÈT�È=��9�l��b@|��� }~�Q����RSD����N8���  '���ap?��P�b!p�b){�B���?�CIpB  X���ذ��C�A�av/ � {��	�o�Q�IB P��8�����P��ԕرD �O���O���A�,�>�Š
�`l�1�	 �٠p��� p` �l`:Ѳ��a�1a�?�ff{O��įV� �P����aa�!��/�?Y)R�a4�(ذ]�Pf����a\c\d^ƃ?333-d����;�x5;��0�;�i;�du;�t�<!�+}�oݯ��b�Sb�P�?fff?��?&���T@��A{#$�@�o[,� ��x�	�&f6�ed�g ���Hd㯸ϣ�����  ���$��H�Z�E�~���&eF��mߺ�i߀��U���y���2���E�0����y�d�� ������������ ?�*�܏r�8�.o�ߺ� ���T�);ڿ Pb��������P��A��T C�=�ϵ��Y}��2������m�C��W�C�= �` Ca��������(!�`�<����bC@_;C9��BA��Q�>V{È�����Y�?uü��
/�S���Q��hQ��A�B=�
�?h�Ä/iP�����W��ÈK��B/
=�����Ɗ=�K��=�J6XK��r#H�Y
H}���A�1�L��jLK����H:��H�K��/0	b�L �2J��8�H��H+UZBu�a?�/^? �?�?�?�?�?�?O�? O9O$O]OHO�OlO�O �O�O�O�O�O�O#__ G_2_k_V_{_�_�_�_ �_�_�_o�_1oo.o goRo�ovo�o�o�o�o �o	�o-Q<u `������� ��;�&�K�q�\���΀�Gϭ���� C�aɏ Ĉ�y���CVF������+b�����yKc�f�� 
E��Ў�T�ٟt�(t��_3�h۟���������N�������3�lC�(�:�H�����T�f��t�.3礁}����k����q'�3�JJ �����گ���4�"�J]P̲Pf��������⟛�ſ���ԻA����/��?�{?�<N�u�  fUh�*� �Ϟ������Ϣ�t�.��R�@��X�bߘ�̆ߨ�)Z�ߺ�  ( 5�	�������B�0�f�t�  �2 E%p"E[[@��N�"B,C��%@ߏ��"����	����?�^������@����%n�n�%T��%��Xc
 ��!3EWi {��������b*[��P�I��v�$MSKCFMAP  ��� ^������pDONREoL  X�[���DEXCFEN�B�
Y�FN�C��JOGOV�LIM�d��d�DKEY��%_PAN�"".DRUN��>#SFSPDTYw�x���SIGN�>�T1MOT���D_CE_GRoP 1���[\���/��?&?��? Q??u?,?j?�?b?�? �?�?O�?)O;O�?_O O�O�OLO�OpO�O�O �O_%__I_ _m__�f_�_O�DQZ_E�DIT�$UTC�OM_CFG 1��Q�_o"o
��Q_ARC_��X��T_MN_M�OD���$�U?AP_CPLFo��NOCHECK {?Q W� ���o�o�o�o' 9K]o������vNO_WAI�T_L�'�W� NT��Q�Q���_7ERR�!2�Q��� �_t�������A*��Ώ�d``OI�}�P�x 4��t��C+���XG���k)�70�������8�?0�4�ӏ��|d�B�PARAMJ��Q����_�����s�� =��345678901�� � ���?�Q�-�]������u���ϯ����������7�ODR�DSPEc�&�OF�FSET_CAR8�PKom�DISz�K��PEN_FILE����!$a�V<`OPT?ION_IO
/=!�аM_PRG %Q%$*	�ά�WORK ��'=� ��Kƪ�P��/����f�(�f�	 ���f�5����M�RG_D?SBL  Q������L�RIEN�TTO* ��C����Z��M�UT_S/IM_DطX+�M�VQ�LCT ��%��R_�$aQ�'�_�PEXh`��b�RA-Thg d�b�r��UP �5� �� ����߼������$��2�#�L6�(L?��	l d'�O�a�s�� ������������ '�9�K�]�o���������H�2>������/ASew�N�< �������@1CUgyH����P�� � � ��  �U�A��  B��PB�����H���  ���U�BJ�p������N��P Ez  E��� E�` EE��;(�����Z�/���  �E��''���@V#���T�AJ(��E!Y!a!)!m!Y!�u)%)!Y!E!�%E!��$�^$A!�	!E!a! �%%	-Y!Y%�-58��Z 99U%E!�D!	$D%%E!Q481X2 91�%�)95�/W#95)%�91m5a!�5/Z7��Z (�8�1�<a1 fEE	�(�Em�4�94X6E9=)%E15�� |O�O�O�O�O�O��O�O__0_B_T]F�S_y_�_�_�Vh������_�[��͔ on�_=oKg�]�]&��'4 � �W%po�oX� Н��g�o�jA�A��c�����o�o$*w���tB�(~ ΐ��r�|�` q�y��$�O��1�-�k�-��3��`��0��P( @EhD�D��q?Q�C�Z7�}��o  ;�	l�D�	u� ���pX��[�2��X �? � �,i�X��ΐH��9H��H��H`��H^yH�R�l���_����	�#�5B#�B C4ӄ�����c�9���
=���� �������cBz���Βa�m� 另b�s�� �q���gd䟒�챏Ǒ�ٖ��o���e	'� �� �I� ��  �q<�=����9�K�E�@a�g�b���������!E������N�㯇  '۰��Ɓ"�B��Ղ��т6��� ~�  ��C�aB��	ŀ~��p=�Bp ��Н����px����D��o޿�o��&�l�#�5�Ю`Q���	 ٠TU�f� U� Q�:����#����?�faf\o�ϩ�;� �p�����F�8� ��?%Y
r��q=�(� BՁPK�fɆ�A�A���?�333��Ł;��x5;��0;��i;�du;�?t�<!��y�������t���r�p?f7ff?x�?&����@��A#	�@�o[�	]� �����uI��wh��� -��ϝ��������� 	���-�?�*�c�u�L� ������4�V�X����EjPf��^ I�m����  �$��W� ������9��/  /��5/G/�z/e/�/`�/�/�/�`�A��$�t�/ C�/"?�(d��>�?��Pn?�/h�?}?��(��W�?{C�@�` CT���?�j4�j0i1A@�I�!���bC�@_;C9�B�A�Q�>�V`.È�����Y�uü��
�?�3��Q���hQ�A��B=�
?h���iOJp��W���ÈK�B/�
=�������=�=K�=�J�6XK�r#H��Y
H}��A��1�=L�j�LK����H:��HK���O�@	bL ��2J��8H���H+UZBu�?F_�OC_|_g_�_ �_�_�_�_�_�_o	o Bo-ofoQo�ouo�o�o �o�o�o�o,P ;`�q���� �����L�7�p� [��������ȏ�ُ ���6�!�Z�E�~�i� {�����؟ß��� ���0�V�A�z�e�G�y����� C�a�/>�� Ĉ��ЯׯOCVF�����üK<G�b0��KH�K�� 
Ep�s�9���z� (�!�_�h���y����a5�N�����T�3lC�8��-¢�9�K���t�.3��}�e�w�k���q'�3�JJ�͑���@��������B5P��	PK�Zgt�ǿ��0�ߕ��߹�����߈���$�{$�3�Z�  fUM����� �����Y��7�%���=�G�}�k���)�Z����  ( 5�� ������'�KY  2 wE%pIFE[@t�N�IFB�!�!� C%��0� T�@į�����*H3 ��Tfx��T�T�a4��T�D9=4H;
 �/ /*/</N/`/r/�/�/��/�/�/�/�/GJ@2���5�I�v�$�PARAM_ME�NU ?����  �DEFPULS���	WAITT�MOUTT;RC�Vg? SHE�LL_WRK.$�CUR_STYLv���<OPT�N�?PTB�?�2C�?R_DECSN_0 <�L	OO-OVOQOcO uO�O�O�O�O�O�O�O�_._)1SSREL?_ID  ��Y��=UUSE_PR_OG %8:%*_�_>SCCRk0ORY�@3�W_HOST !8:!�T�_�ZAT\Ю_ c�_�Qc|<o�[_TIMEi2�OV�U)0GDEB�UGMP8;>SGIN?P_FLMS`�gn�hTR�o�gPGA��` �lC�kCH��o�hTYPE5<A)_#_Y�}� �������� 1�Z�U�g�y������� ������	�2�-�?� Q�z�u�������ϟ��
��eWORD �?	8;
 	�PR�`U�MAI�@��SU�1E�T1E#`U��	�4R��COLS�n���vT�RACECTL �1���B1 ]W ] �W �d�ެ��DT Q����РD �� ;�* eZ �d� � �6��6��`6�ۡ7�T�6�4�2�:�UB�4�	4�
4�U4�2�:�B�4�4�(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v�������0*<�\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhzP ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� �0�B�T�f�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼� �������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�?��?I�$PGTR�ACELEN  �A  ���@�$F_U�P ����2SA[@?AT@$A_CFG �SES=CAT@��D��D�O�G6@�OhBD�EFSPD ��sLA6@�$@H�_CONFIG s�SE;C @�@dT�3B �AQP�D�A1Q@��$@INk@TRL' �sM�A8�EFQ�PE�E�W��SA�DQ�ILID�lC�sM	�TGRPW 1�Yb@lA�C%  ��l��AA��;H�N���R���A!PDg	� a3C	\T�Ai)iQP� �	 �O4VGgCo #´|c^oGkB`�a��opo�o�o�o�o�b?"�Bz�o7�I~3 <}�<�oN�J�� ���f�)��9��_�J�`z����@
 t���d�ŏ�֏��� 3��W�B�{�f�x������՟�����J)@)�
V7.10b�eta1�F �@�@�OA&ff�Q2�CPkC�`�D�Dk`�[�C�T��@ DĠ Dr� �Q�BH�`�L��PC5zR A?�  ��#CCx����b��P!P���A����Ap�B<�b!PA1�������
�?L��?33�3A@��"��Ff�f.��b�w:�7���AeC�QKNOW_M  �E|{F�TSV �Z(R�C������ʿ ��ٿ�$�A!m�SuM�S�[ �B��	�E���PϏ�̓E`��2�E�@�2�������� VL�MR�S�Y�T�j	���AC5����e@��Rۚ]ST�Q1 1=�SK
 4�U��A�¨߰E��*��߽� ������J�)�;�M� _�q��������� ���F�%�7�|��Ep��2{���A�<�����P3���������p�4��+p�5 HZl~p�6����p�7� $�p�8ASewp�M�AD0F [Fp�O�VLD  SK��ϼOr�PARNU�M  /�O//T�_SCH� [E
�}'F!�)=C�%UPD�F/X)�/3Tp�_CM�P_O�0@T@@'�{E�$ER_CHK�5yH!6
?;RS8�]��Q_MO�o?�5_k?��_RES_GzФ~ݍ��?�O O�?%OO*O[ONOO rO�O�O�O�O�O�O��3���<�?_�5�� (_G_L_�3G g_�_�_ �3� �_�_�_�3� �_ o	o�3@$oCoHo�3��co�o�o�2V 1�~կ1e�@c?���2THR_IN�R�0�!7³5d�fM�ASS ZwM�N5sMON_QUEUE �~�Xf��0�� �4N0�UH1NEv6;�pENqD�q�?�yEXE���u� BE�p��sO�PTIO�w�;�pP�ROGRAM %hz%�p�ol/�r?TASK_I��~OCFG �hx/\���DATAR�]���@��2�� ���#�5�G��k�}� ������^�ן����^��INFORé܍�wtȟe�w������� ��ѯ�����+�=� O�a�s���������Ϳ4(�4��܌ �I��6� K_�����T��ENB� ͻ1>�h��I��G��2��? P(O�ҡώ�� �����_EDIT �����ߋ�WERFL��x�cm�RGADJ7 �8�AС�iԁ?�0t�
qLֈq����5�?��!��<@��*�%����@�#ߊ��2����F�	Hpl�G|�b��>��A�dw�t$I�*X�=/Z� **:c�0 V�h���Ǟ���B������������� ������b���L�B� T���x���������: ����$,�Pb ������� ~(:h^p� �����V/ // @/6/H/�/l/~/�/�/ �/.?�/�/?? ?�? D?V?�?z?�?O�?�? �?�?�?rOO.O\ORO dO�O�O�O�O�O�OJ_ �O_4_*_<_�_`_r_ �_�_�_"o�_�_ooo�f	���o�p�o�o �dJ��oL��o#�oG�Y��PREF �����p�p
L�I�ORITY����>P�MPDSP�>�ƴwUTz�4�K�OD�UCTw�8��\�OG�_TG�;�|����rTOEN�T 1��� (�!AF_INE��pp�{�!tc�p{���!ud���ˎ!icmX�����rXY�Ӵ��;��q)� p�/�A��p�)�j�M�Y� ��}��������ן� ��8�J�1�n�U�����	*�s�Ӷ}}�����^,�>��jfp�!/z�֯K�,�������A��,  � �p�������ʿ�u"��ut�}�sF�P�PO�RT_NUM�s��p�P�_CARTREP�p��|��SKSTA�w nK�LGSm���������pUnothingϿ�������c{t�TEMP �����ke��_�a_seiban 0C�,S�y�dߝ߈� �߬�����	����?� *�c�N��r���� �������)��M�8� q�\�n����������� ����#I4mX �|�������3��VERSI��p �d disabled>SAVE ���	2600H7K21:&�!;�0��̏� 	(�r$moN+E/`�eb/�/�/�/�/�*z,�?� %`���_-� 1���E0�b8e�O?a?4gnpURGE_ENB3��v�u�WF�0DO�v��v�Wi��4�q*�WRU�P_DELAY ��CΡ5R_HOT %�f�q:�.O��5R_NORMA�LH
�OrOAGSE�MIQOwO�OlqQS�KIP-3���>3x $�O _1_C_]&o t_b_�_�_�_�_�_�_ �_o(o:o o^oLo�o �o�olo�o�o�o  $�oH6X~�� h��������D�2�h�z�����$�RBTIF�4G�R�CVTMOU\�v����DCR-3}��I �Q�=���1D�a��Ab�S<8@��3�.?�[��-�Ģ�lQU�?����\�_�X�T_;�x5;���0;�i;��du;�t�<!���h��R���̝ �����&�8�J�\��n����������RD�IO_TYPE � 4=��¯EFP�OS1 1�C�
 x/:�H2��b�M� ��/��E�οi�˿� ��(�ÿL��pς�� /�i��ϵ��ω�߭� 6���3�l�ߐ�+ߴ� O����߅ߗ���2�� V���z���9���� o�������@�R������9��������OS/2 1��;+�u����-��Q���3 1�����G��|�gS4 1�~����ZE~�S5 1�%7q���/�S6 1Ũ��/�/o/�/>&/S7 1�=/O/�a/�/??=?�/S8 1��/�/�/0?�?��?�?P?SMASK 1�߯ )�OFN�7XNOܯFUO<_C�MOTE����X4uA_CFG ��|M�1\A�PL_�RANGxA���AO�WER ����@�FSM_DRY�PRG %�%�y?!_�ETART ���N/ZUME_�PRO�O_�_X4_�EXEC_ENB�  ����GSP�DdP�P�X���VTD�B�_�ZRM�_�XI�A_OPTION�φ����pAINGoVERS.a��z_�)I_AIoRPUR�@ @O\�o�=MT_�0T�@�zO��OBOT__ISOLC=N�F��1�a�eNAME�Rl�bo�:OB_O�RD_NUM ?��H�aH�721  V1;wLqr�qrV0.qr��sps�u�\@��PC_TIM�Ė��x��S23�2�B1����aL�TEACH PENDAND��1\H���x?c�Ma�intenanc�e ConsV2��#�"�_�No Use��N��r����������С�rNPQO>P�r\A<e�qoCH_LgP�|N�w�	<��!U�D1:b�	�R�0VgAILRq2e��u�pASR  ��:a�B�R_INoTVAL1f��I��+n��V_DAT�A_GRP 2�X��qs0DҐP�? `��?��o�������� կï�����-�/� A�w�e���������� ѿ���=�+�a�O� ��sϕϗϩ������ ��'��K�9�[߁�o� �ߓ��߷��������� �G�5�k�Y��}�� �����������1�� U�C�e�g�y������� ������	+Q?�uDA�$SAF_DO_PULS�p�E@�C�� CANd�r1f�vpSC�@��-�-�}��QV0D�D�qL�L�+AV2 y�'9K] o��������ڈ��2$($Md($C!u�1#
) @�Co/�/�/ȥ.W)k/ M��$_�_ @݃T:`��/??&?39T D��3?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O֏��i%�O�O�O܉x�!L� �;�o݄��p�M
�t��Dipp�L��J?� � ��jL� ��j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt ���������(�:����/c�u� ��������Ϗ��B� %�1�C�U�g�y���@������Ƒ��0R MS�EW]�$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ�����M���*� <�N�`�r߄ߖߨ�� ��������&�8�J� \�ǟ���������� ��������,�>�P� b�p������������� ��%7I[m ��������!3EWit�OB3t���� �////A/S/e/w/@�/�/�/�/�/�*���/?6��\R�?�M	1234�5678XRh!?B!̺����?�?�?�? �?�?�?OOA�>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ o]-O�_�_�_�_�_�_ �_o"o4oFoXojo|op�o�o�oq_BH�o �o�o!3EWi {�������<�v[;�j�A� S�e�w���������я �����+�=�O�a�xYD�k�������ɟ ۟����#�5�G�Y� k�}�������v_ׯ� ����1�C�U�g�y� ��������ӿ���	� ȯ-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�σߕߧ߹� ��������%�7�I�[�m�����v6����z��!�3��O:Cz  Aоz   �@�2��v0� @�
~���  	�r�������������ph�u�����K] o������� �#5GYk} ��0����/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-?�G�������*@  <�X4t��$SCR_�GRP 1�-�� -�� t� �t� �E5	 �1��2�2�4�� W1G3�;97�7�?�?O�C��|�BD�` D��3NGK�)R-200�0iC/165F 567890���E��RC65� �@�
123I4�E�6t�A�����C�1F�1�3�1�)�1A�:�1�I	���?_Q_c_u_�_���H��0 T�7�2�_�?�_�_o�6�t��_Lo�_poB8�boK�h�@�UO��q  NM�1B����B�  B�33Bƿ`�e�b�cr�1Ag��o  @t���e�1@>@	  ?	�w�bH�`2�j�1F@ F�`\r d[o�s���� ���*��9�a�a)r`U�@�R�d�v�B��� �ʏ���ُ���� H�3�l�W���{���@Ě2C�?���7����9�t�!q@"p>�1?�S�r�`y��`ȏ��G�L�3��ϯ�A>G�1��"oeI��)�t� �<�N�\�*�q�}���.^� P��(�����ӿ�g1EL_DE�FAULT  ~�D��t����HOTSTR�� ��MIPOWERFL  K�x���?�WFDO�� S�RVENT? 1����P0�� L!DUM�_EIP翬��j�!AF_INEx��ϵ!FT�ϒ�����!�_B� ���i�!RP?C_MAINj�L�q�Xߵ�|�VIS���Kٻ���!TP&��PU�߳�d��M��!
PMON_POROXYN��e<��g��f����!�RDM_SRV����g��1�!RȻDM���h �}�!
�~�M���il���!?RLSYN�@�����8��!R3OS��<�4a�!
CE�MTC�OMb��kP�!=	vCONS����l��!vWA'SRC ���m�E;!vUSBF��n4�0ߵ��� �/�'/�K//o/��RVICE_K�L ?%�� (�%SVCPRG�\��+�%2�/�/� 3��/�/� 4??� 5�6?;?� 6^?c?� 7@�?�?� �D�?�,9�?�;�$H�O�!�/+O �!�/SO�! ?{O�!(? �O�!P?�O�!x?�O�! �?_�!�?C_�!�?k_ �!O�_�!AO�_�!iO �_�!�Oo�!�O3o�! �O[o�!	_�o�!1_�o �!Y_�o�!�_�o�!�_ {/�"� �/� F�E1 �������� 
�C�U�@�y�d����� �����Џ����?� *�c�N���r������� �̟��)��M�8� _���n�����˯��� گ�%��I�4�m�X� ��|�����ǿ�ֿ���*_DEV ~���MC:��H'�GRP 2�ׇ�+p� bx 	� 
 ,y�ϒ�+r~ϻϢ��� �������9� �]�o� Vߓ�z߷��߰����� �#�z�G���k�}�d� ������������� ��U�<�y�`����� ����*���	��- QcJ�n��� ���;"_ FX������� �/�/I/0/m/T/ �/�/�/�/�/�/�/�/ !??E?W?�{?2?�? �?�?�?�?�?O�?/O OSO:OLO�OpO�O�O �O�O�O_^?�O=_�O a_H_�_�_~_�_�_�_ �_�_o�_9oKo2ooo Vo�ozo�o�o _�o�o �o#
G.@}d �������� 1��U�<�y����o�� f�ӏ�̏	���-�?� &�c�J���n������� �ȟ����;���0� q�(���|���˯��� ֯�%��I�0�m�� f�����ǿ������R�d ��	�4���X�C�|�gϠϯ�%�x����R������ ���������+��O� =�s߁��Ϧ���i��� �������	��Q�� x��A�������� ���Y��P���)��� q�����������1� U���I��Ym� ��	�-�! E3U{i��� ���//A/// Q/w/��/�g/�/�/ �/�/??=?/d?v? -?O?)?�?�?�?�?�? OW?<O{?OoO]OO �O�O�O�O�O/O_SO �OG_5_k_Y_{_}_�_ �__�_+_�_ooCo 1ogoUowo�_�_�oo �o�o�o	?-c �o��oS�O�� ���;�}b��+� ��������ɏ�ݏ� U�:�y��m�[���� ����ş�-��Q�۟ E�3�i�W���{���� دꯡ�ï���A�/� e�S���˯���y�� ѿ����=�+�aϣ� ��ǿQϻϩ������� ���9�{�`ߟ�)ߓ� �߷ߥ�������A�g� 8�w��k�Y��}�� �������=���1��� A�g�U���y������� ���	��-=c Q������w�� �)9_�� �O����/� %/gL/^//7/// �/�/�/�/�/?/$?c/ �/W?E?g?i?{?�?�? �??�?;?�?/OOSO AOcOeOwO�O�?�OO �O_�O+__O_=___ �O�O�_�O�_�_�_o �_'ooKo�_ro�_;o �o7o�o�o�o�o�o# eoJ�o}k�� ����="�a� U�C�y�g�������ӏ ���9�Ï-��Q�?� u�c���ۏ��ҟ���� ���)��M�;�q��� ��ןa�˯��ۯݯ� %��I���p���9��� ��ǿ��׿ٿ�!�c� Hχ��{�iϟύ��� ����)�O� �_���S� A�w�eߛ߉߿���� %߯���)�O�=�s� a���߾��߇����� ��%�K�9�o���� ��_����������� !G��n��7�� ����O4F ��g���� �'/K�?/-/O/ Q/c/�/�/�/��/#/ �/??;?)?K?M?_? �?�/�?�/�?�?�?O O7O%OGO�?�?�O�? mO�O�O�O�O_�O3_ uOZ_�O#_�__�_�_ �_�_�_oM_2oq_�_ eoSo�owo�o�o�o�o %o
Io�o=+aO �s���o�!� ��9�'�]�K���� ����q���m�ۏ��� 5�#�Y�������I��� ��ßşן���1�s� X���!���y������� ��ӯ	�K�0�o���c� Q���u��������7� �G��;�)�_�Mσ� qϧ����ϗ�ߓ� �7�%�[�I���Ϧ� ��o����������3� !�W��~��G��� ��������	�/�q�V� �����w��������� ��7�.����O �s����3 �'79K�o ������#/ /3/5/G/}/��/� m/�/�/�/�/??/? �/�/|?�/U?�?�?�? �?�?�?O]?BO�?O uOO�O�O�O�O�O�O 5O_YO�OM_;_q___ �_�_�_�__�_1_�_ %ooIo7omo[o}o�o �_�o	o�o�o�o! E3i�o��Y{ U�����A�� h��1����������� ����[�@��	�s� a������������3� �W��K�9�o�]��� ��������/�ɯ#� �G�5�k�Y���ѯ�� ����{�����C� 1�gϩ���ͿW��ϯ� �������	�?߁�f� ��/ߙ߇߽߫����� ���Y�>�}��q�_� ���������� ������7�m�[���� ����������� !3iW������ }���/ e���U��� �/�/m�d/� =/�/�/�/�/�/�/? E/*?i/�/]?�/m?�? �?�?�?�??OA?�? 5O#OYOGOiO�O}O�O �?�OO�O_�O1__ U_C_e_�_�O�_�O{_ �_�_	o�_-ooQo�_ xo�oAoco=o�o�o�o �o)koP�o� q������C (�g�[�I��m��� ����ُ� �?�ɏ3� !�W�E�{�i����� ؟������/��S� A�w�����ݟg�ѯc� ����+��O���v� ��?�����Ϳ��ݿ� �'�i�Nύ�ρ�o� �ϓ��Ϸ�����A�&� e���Y�G�}�kߡߏ� ������ߵ��߱�� U�C�y�g����������$SERV_MAIL  ������OUTP�UT���RoV 2؍�  �� (����_���S�AVE���TOP�10 2�9� d 	�������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/����YP|���FZN_CFG ڍ�'��j��!?GRP 2��'&�� ,B   A�=0��D;� B�>0�  B4���RB21l�HELL�"܍�$�L��M�7�?�;%RSR�?�?�?O�?%O OIO4OmOXOjO�O�O��O�O�O�O_!_3^�  �R3_a_Xs_AR_ ��{_L�R�P�xWIR2���d�\�]�Rh6HK ;1�v; �_o "ooFooojo|o�o�o �o�o�o�o�oG�BTfb<OMM ��v?�g2FTOV_ENB��A�$���ROW_REG_�UI���IMIO/FWDL�pߥ~@5^�WAIT�r�Y��8���v@�0�T�IM�u��j�V�A��A��_UNI�T�s��$�LC�pT�RY�w$���M�ON_ALIAS� ?e�yH�he ��%�7�I�[�i���� ����m����
�� .�ٟR�d�v�����E� ��Я������*�<� N�`��q�������̿ w����&�8��\� nπϒϤ�O������� ��߻�4�F�X�j�� �ߠ߲����߁���� �0�B���f�x��� ��Y����������� >�P�b�t�������� ������(:L ��p����c� � �6HZl ~)������ / /2/D/V//z/�/ �/�/[/�/�/�/
?? �/@?R?d?v?�?3?�? �?�?�?�?�?O*O<O NO`OO�O�O�O�OeO �O�O__&_�OJ_\_ n_�_�_=_�_�_�_�_ �_�_"o4oFoXooio �o�o�o�ooo�o�o 0�oTfx�� G������,� >�P�b���������� Ώy����(�:����$SMON_D�EFPRO ����c�� *SYS�TEM*M�REC�ALL ?}c�� ( �}-co�py frs:*�.dt virt�:\temp\=�>192.168�.56.1:10496 ɕ؟�����}xyzrate 61��Αß�՟f�x����8��o�rderfil.�da��mpbac�k��U����� }]/��mdb��*���ʯӯd�v����3x��:\,���>�N�W�P�����4��a�� ��I�ؿi�{ύϠ��� ;�V���������B� ��e�w߉ߜ�/�A�ҿ �����ϫ߽�P�a� s��Ϫ�3������� ��(���L�]�o��� �ߦ�9����������$��H���k}
#� .@R����#�D�8220� ��dv��  .@R��/�,�16���e/w/�/ ���7�8'�/�/�/� $��/7(�/d?v?�?�� ,?�<#W?�?�?O �?�?��?iO{O�O�/ �/;?V?�O�O_?�O B?�Oe_w_�_�?/OAO �?�_�_oO�_�_PO aoso�o�O�O3_�O�o �o_(_�oL_]o ��_�_9o�_��� o$o�Ho�k�}�� �4�F�X����� ��7188�ҏc��u����etpdiosc 0-�8 ?��Q������ftp?conn 0��� ̟]�o����k7�o�oB��8�������.#���6�үc�u����e2 ���2�V����Ϟz +���9�׿h�zόϟ� ��:�U�����
�����A���d�v߈ߚc�$�SNPX_ASG 2��������  �Z�%�����  ?����PARAM ����� ��	��P�d�`���*����OFT�_KB_CFG � �c�՞�OPI�N_SIM  
��%��������RVQSTP_DSBk�%�����SR ���� & CONgROD��/����TOP_ON_ERR  /�W�L�PTN ����AH�RI�NG_PRMV� ���VCNT_G�P 2��'��x 	�����`�� ���$��VD��RP 1���(��� _q������ �%7I[m �������� /!/3/Z/W/i/{/�/ �/�/�/�/�/�/ ?? /?A?S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_r_ o_�_�_�_�_�_�_�_ �_o8o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c����������� Ϗ����)�P�M� _�q���������˟ݟ ���%�7�I�[�m� �������ܯٯ�����!�3�=PRG_�COUNTL��8�[�_�ENB��Z��M��N䑿_UPD� 1�� T  
H���ۿ���(� #�5�G�p�k�}Ϗϸ� ������ �����H� C�U�gߐߋߝ߯��� ������ ��-�?�h� c�u��������� ����@�;�M�_��� �������������� %7`[m� ������8 3EW�{��� ���/////X/ S/e/w/�/�/�/�/�/ �/�/?0?+?=?O?x?�s?�?Q�_INFOg 1�ɹ�� �F���?�?�?O�9����hA��>�>�O�3A���A��3�9�z��Ң�����P�YSDOEBUGi�ʰ�0�d��z@SP_PA�SSi�B?�KL�OG �ɵʴ��0>H�?  �����1UD1�:\�D�>�B_MPAC�Mɵ:_L_ɱ�A�j_ ɱVSAV ���MA�A�B�5� XSVnKTEM�_TIME 1��G�� 0�0̢�4�lX�Z�4��T1SVGUNSİ�j�'���`AS�K_OPTION�i�ɵ����?a_D�I�@��[eBC2_?GRP 2�ɹ�U��o�0@�  C���cP��`CFG ��km�V�f`
OB-Rxc �������� �>�)�b�M���q��� ������ˏ��(�� L�7�p����4m��� n�ϟ�\�����;� &�_�q^�QdT����� ��ѯ�������)� +�=�s�a��������� ߿Ϳ���9�'�]� Kρ�oϑϓϥ����� ������1�C���g� U�wߝߋ������߳� 	���-��Q�?�a�c� u����������� �'�M�;�q�_����� ����������7 ��Oa��!� ����!3E iW�{���� �/�///S/A/w/ e/�/�/�/�/�/�/�/ ??)?+?=?s?a?�? M�?�?�?�?O�?'O O7O]OKO�O�O�OsO �O�O�O�O_�O!_#_ 5_k_Y_�_}_�_�_�_ �_�_o�_1ooUoCo yogo�o�o�o�o�o�o �?!?Qc�o� u������� )��M�;�q�_����� ��ˏ���ݏ��7� %�G�m�[�������� ٟǟ����3�!�W� o�������ïA�� կ����A�S�e�3� ��w�����ѿ���� ��+��O�=�s�aϗ� �ϧ��ϻ������� 9�'�I�K�]ߓ߁߷� m��������#��G� 5�W�}�k������ �������1��A�C� U���y����������� ��-Q?uc ������� ��/A_q�������/� ��$TBCSG_G�RP 2���  � � 
 ?�  J/\/F/�/j/�/�/��/�/�/�/;#"*#�~1,d0?1�?!	 HD� 6s33[2�\5O1B�!x?�9�D)�6L�͞�1>���g6�0CqF�?�?�8fff�1�>��!OICj��6�1H4B�GC{OO)H��02|A�]0@HDO_O�)H�1�8CFr�O�M@  �. XU&_�O_Q_�n_9_K_�_�_�[?���0�Sp �	V�3.00�R	rwc65�S	*`��T"o�V|A�0 8 `�Y G`mHoW  � �%@�_X�o�c#!J2*#�1-��o�hCFG ���;!C!�j��B"]b�l|�BPz�Pva �������� �<�'�`�K���o��� ����ޏɏ��&�� J�5�n�Y�k�����ȟ ������\	��-� ן`�K�p��������� ޯɯ��&�8��\� G���k�����!/ۿ �����5�#�Y�G� }�kϡϏϱ������� ����C�1�S�U�g� �ߋ��߯�����	��� �?�-�c�Q���Y ����m������)�� M�;�q�_��������� ��������%I[ m9����� ��!E3iW �{�����/ �///?/A/S/�/w/ �/�/�/�/�/�/?+? ��C?U?g??�?�?�? �?�?�?�?OO9OKO ]OoO-O�O�O�O�O�O �O�O_�O!_G_5_k_ Y_�_}_�_�_�_�_�_ o�_1ooUoCoyogo �o�o�o�o�o�o�o 	+-?uc�� ��y?����;� )�_�M���q������� ݏ�����7�%�[� I��������o�ٟǟ ����3�!�W�E�{� i���������ï��� ��A�/�e�S�u��� �������ѿ���� �+�a��yϋϝ�G� �ϻ������'��K� 9�o߁ߓߥ�c��߷� ������#�5�G��� }�k���������� ����C�1�g�U��� y�����������	�� -Q?a�u� ������/ ���q_���� ���/%/7/�/ m/[/�//�/�/�/�/ �/?�/?!?3?i?W? �?{?�?�?�?�?�?O �?/OOSOAOwOeO�O �O�O�O�O�O�O__ =_+_M_s_a_�_C �_�_}_�_�_o9o'o ]oKo�ooo�o�o�o�o �o�o�o#Yk }�I����� ����U�C�y�g� ��������я���� 	�?�-�c�Q�s�u��� �����ϟ��)�;� �_S�e�w�!�����˯ ��ۯݯ�%��I�[� m��=�����ǿ����վ  �� ��)���$TB�JOP_GRP �2�ݵ��  ?��	�A�H��O���� ����pXd� ����� � �=,� @�`�	 �D ���CaD����`���fff��>���H�ϻ�L���	�<!a���>����=�B�  �Bp��8�C�D)��U�CQp�D;�S�Ι��y����v� ?�������\<���U��[��%�CV+��/�<��S�D5mi�{����ع�<�����z�>\>��33C�  CA8��`�K�j��u�b�����z�;�9b�B�E�>�}׵ҳ� C�V����s����&��ǌ��;��6��%�]�?D&� C���������
Ѷ� ?s�33����<Z;u����ff�ҴK�� ����U�)C-_ i�u����� �*IcMH�����Ƙ����	V3.00f��rc65e�*� e��/ ' �F�  F�� �F� F�  �G� GX �G'� G;� �GR� Gj` �G�� G�| �G� G�� �G�8 G�� �G�< H� ?H� H��2 �Ez  E�@ _E�� EB F� �FR FZ F�� F� F�P<"G � GpL#�?h GV� G�nH G�� G��� G�( =u=+�(�$`Q�?2��3?�  ���M?[:A��*S�YSTEM
!V8.30218 �3�8/1/2017� A y  �p7M�TP_TH�R_TABLE   $ $�1�ENB��$DI�_NO��$DO��4  ��1CF�G_T  0��0MAX_IO_�SCAN�2MIN��2_TI�2DME�\��0@�0 � � $COM�MENT ]$CVAL	CT�0�PT_IDX���EBL�0NUMQBE�NDIJfAZITID�]B $DUM�MY13��$P�S_OVERFL[OW�$�F�0wFLA�0YPE�2��BNC$GLB_�TM�7�EF@�1�0O�RQCTRL�1��$DEBUG��CRP�@2@  �$SBR_PA�M21_VP �T$SV_ERR�_MODU4SCL|�@RACTIO�2��0GL_VIEW��0 4 $�PA$YtRZtRW�SPtR�A$CA�@A�1�_SUeU� �0N�P3@$�GIF3@}$eQ �lP_S�PiQ L�pP�VI<P�PF�RE��VNEARPLA�N�A$F	iDI�STANCb�1J�OG_RADiQ�@$JOINT�SP尤TMSE]TiQ  �WE�UACONS2@B�R�ONFiQ	� �$MOU1A`��$LOCK_FOyL�A�2BGLV@C�GL�hTEST_sXM@@raEMPE`�,R�b�B`�$U1S;AfPH`2P�S:�a�bMP_�`�a=QCENEdRr� $KARE�@M>�3TPDRAhP;t>2aVECLE�32dkIU�aqHE�`�TOOLH`�0qsV�I{sRESpIS3�2�y64�3ACH4X`�`~qONLE�D�29�B�pI�1 � @$RAIL__BOXEHaPoROBO�d?�Q?HOWWAR�0�r<�@�qROLM�B�A�C �SK�r�@�07O_F9�!��St�qiQ
>o �RVp�OCiQ_�SLO�GaK��VOUZb�R�eAELEC�TE<P`�$PI=P�fNODE�r�r��qIN�q2^��pCORDED�`�`}��0P9P@  wD �@OBAU`TA�a����C�@��p�P�q0��ADRAܥ0F@TCHup 7 ,�0EN�2�1A�a_�Tl�Z@�BޣRVWVA!A� � ApeR�5P�REV_RT�1�$EDIT��VS�HWR9�S@	UАI�S`yQ$IND�0@1QB蓗q$HEAD�5@ ��p5@溒KEyQ�@CPS�PD�JMP�L��5�0RACE�4U�a�It0S�?CHANNEzp��	WTICK{s�1M�`A�0@�HN�A�D0^�]D�`CG�P8���v�0STYf��q�LO�A�3B���jP� t 
��Gr�%�$���T=PS�!$UNIGa5A�E��0�FPORT��SCQU5ptR���B��TERCJ@���T=SG� �PPL6�$�DE��$`Thqb�0OK@>CV�IZ�D4�Q�E�APR�A�Ͳ�1��PU}aݵ_�DObk�XSV`KN�6AXI��7�qgUR_s�E$T�p���*��0FREQ_,hp<�ET=�P�b�OPARA`@.P
@�:[���ATHr�3@a�D�s�s�0 �2�SR_Q�0l8}��@�1TRQIc���$`�@��BRup��VyE@@��NOLD��AAp7a��x@�A��AV_MG����¨/���/�D)�D;�D�M�J_ACC.�C��<�CM��0CYC0M@3@��M@_E������٘@NbSSC��@  hPD1S���1�@SP�0*�AT:����@��i��B�ADDRES{sB���SHIF}b�a_W2CH�@&�I�@�|��TV�bI�2�]��h>��C�
�j
p00����0 \���������웱�@��C�nӞ�aºꯆ:R���TXSCREE���0�TINAWS�P;��T�1>�>�jP TQ�7P�B� 6QP��
��
���RROR_"a�@�؁�E�UEG� ����U��@SXQ�R�SM�� �UNEX0g��6��0S_�S@��	0��>�C�b���o� 26�UE���2GRUͰGMTN_FLQ��#POHgBBL�_�pWg@�0 �����O�Q�LE�n���pTO`C�RwIGH�BRDIT�d�CKGRg@�T�EX,���WIDTH�sݐB�A�A{q���I_/@H��  8 $LCT_ �|�Y0@RyP@�b�s�w�B��GOu�J�0D0TW� U� r�R�b�LUM�!�^�ERV��]PFQP`>��1'@r�/GEUR�cF\��QM)��LP�Z�Ed��)'�$(�$(�p�#)5!+6!+7!+8 "b�>CȰ`��F�q��aS�@EU{SReT  <���/@U�R��RFOC\hq�PPRIz�m�@�?A� TRIP�qOm�UN�0�4!�P ��0�5�7��b;��5� "T� ̱G �T7���}�O2OSNAd6RA���;3wq�1#n_�S�^�2��$���aU!"A$�?�?p+"��;3OFF�`� P%O��3O@ G1#PD,D$P�GUN#K`S�B�_SUBBPk SRT�0��&��"avp欳OR�p�ERAU���DT�Ib��VC�C��H�' ��C?36MFB1���PPG?�( (\b`�STE�Qʀ�9PWTѠPE���G�Xd) ����JMOcVE��{Q6RAN4`�?[�3DV�S6RLIM_X�3qV�3qV\XvQ�k\:V1�IP�2V	F��C砽@��G�*��IB�P,�S� _�`�p�b���@/ (0GB�� �"P�@��pr+x# �r �,�tRn�@��s C@TeDRI�PSfQV!�wdԐ���D�$MY_UBY�$\d�;QA�S��q�h�q�bP_S��ף�bL�BMkQ�$j�DEYg�EX�� ���BUM_MUb6�X�D<q US��?��;VGo�PACI�TP�<Uyr�3yr0kSyr:;qREnrጋ1l�9cyr�@,^�BTARGPP�Ⱦp�R<aR{0�@- !d��;cB	:r���R�DSWqp�Sn�$:s˰O�!d�Av�3�
��E��U�p0m���V:cHK�.��K�`AQ��0���?SEA�����WOR�@3��uMwRCVr/ ��UO��M�@C�	Â8C�sÂREF�� ̆��gRj�
�� Ȋ��ي��=�̆r�_RC��s�����@���☩b������to0 �Т�;��� �e�OU���r��\c(`+�u��2��<����̰� -=���f�K��SUL3a.�C�7Po/+p�NT �a��]��ag��g��!g�&�L�c���c�������!�@T��s�1����o@AP_H�UR�ۥSA>SCM�P��F�����_�&�R�T������X�.���VGFS�E2/d �M� � Y0UF_�����J��RO� ����W,rUR�GR�mq�AI���D_V_h[D�@�zY��3�WIN.rH���X-V
A�RqR�P�WEw�w�q|c6v�,q��RvLOiPtc��PMc��3t +�=�PA' =�CACH6����ŵ�,pP����K�ۓC�QIo�FR"�T� $֭�$HO�@�R��`�rc ��[�֘p��ڔ��VP�r����_SZ�3p���6����12�� ��]p�؆P��WA�3�MP��aIMG�x���AD�qI�MREٔ6�_SI�Z�P��!po�6vA�SYNBUF6vV�RTDh�t�F�OLE_2D�T��t�J�0C0aUs��QP��X�ECCU�xVE�M�p����#�VIR9C��VTP������G�p��t��LA@�s�!���Mco4��};�CKLASQCq	��ђ�@5  �AH�� @&B�T$��$`��6 |F@o���Xñ�T�o�?a��"¨uI���r/��`BGf� VEJ�`PK|p`1���֖K�MHO+�>�R7 � }F�x��ESLOW}w�]RO>SACCE0*@-�=�xVR:��11�yrAD�/0r�PA��&�D�1��M_Ba�81��J�MP���A8y�b�$SSC6u��M��$C��@92��S8�ƹN/�PLEX��:# T〲C�Q��6��FLD?1DEZ�F�IQ rO�qty�� K�P2��;�� ϱPV多�MV_PIZ��G�BP0��`а�FIQ�PZ�$��������GA%p�LO9O0Tp�JCBT*����� ��ړPLAN�R&�L�F���cDV�'M�p���U�$�S�P.q�%�!�% #�㱶C4G�����RKE�1�VAN�C]K�A0p <R�@�?�?Q3A�a =�?q??T0�9����r> hܰ�	��!K9�fA2b<X@̠SOUe�ݒA��
O����SK(�M�VI=E�p2= S0:�|R? <{@X��^�`UMMY����jRe��D����A�CU�`b�U�@@� $�@TIT 1�$PR8�UOP�T�VSHIF<ʀ�A`�a����D�0����$�_R$�UړQ.qZ�U �s�ot�Qav�Q5rfSTG@cVSCO��vQCNT���3� }w �RlW�RzV�R�W�R�XPLo^opjjA2��51qD>a�0� �pSMO��B%TC�YJ�@1u���_����@C%�Gi�LIx� '��XVR�D�DY�@T��oZABCP�E�r�b���
�ZIP��EF%��LV��L�����bMPCF��eGy�$p	�~rDMY_LN$@pAr8��dH ����g��>�MCMİC>��CART_Xq��P�1 $JvsptD��|r�r�w��8�u���UXW�puUXEUL�x�q�u�t�u�q�q�y�q�v<�b�eI Hk�dԬ��Y�`D�� �J 8o�	V�EI3GH��H?("��fr��ĔK �= X�C���`$B&�K��b�1_�B��LgRV� qF�`��COVC؀�qrfq9��@}�e�
h����7�D�TRȰr	�V�1�SPH� �ǑL !�S�i�{�����ST�S  ���������� v�<�ѐNa1� ���� ��������������������������	���a��(������������8��( ��RDI������ğ֟����t�O|���������ί���Sz��� >����� ſ׿�����1�C� U�g�yϋϝϯ����� �����v�}���8�!� 3�E�W���'�9�K��]���� ��U��U��� ��8( ��� ���@A�v�^`BF_TAT��ի���I�V>0�n�J�_�I�R 1=&� 8����d%к� ��C�  �� �����������"�4� F�X�j�|��������� ����1gBTjx������р����0B QI�ZlJ�� �������/"/ 4/F/X/FҒ�t/�/b*@���/�/��bv�@`��v�MI_CHANU� `� #3�dV�`哑&0ET>�A�D ?��y0�m��/�/�?�?�d0�RLPs�!&�!��4�?�<SNMAS�Kn8��1255.4E0�33OEOWOտOOLOFS^Q � �%X9ORQC?TRL &�V�m��O��T�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo(l`�OKo:ooo��PE�p�TAIL8�JPGL�_CONFIG �	�ᄀ/�cell/$CID$/grp1so@�o�o1�#��? \n����E� ���"�4��X�j� |�������A�S���� ��0�B�яf�x��� ������O������ ,�>�͟ߟt���������ίB�}c���(��:�L�^���`o��e�� b���Ϳ߿���\� 9�K�]�oρϓ�"Ϸ� ���������#߲�G� Y�k�}ߏߡ�0����� �������C�U�g� y����>������� 	��-���Q�c�u��� ����:������� );��_q��� �H��%7 �[m�����]`�User� View �i}�}1234567890�
//./@/`R/Z$� �cz/���2�W�/�/�/�/??u/�/�3�/d?v?��?�?�?�??�?�.4 S?O*O<ONO`OrO�?�O�.5O�O�O�O_ _&_�OG_�.6�O�_ �_�_�_�_�_9_�_�.7o_4oFoXojo|o�o�_�o�.8#o�o�o�0B�ocir �lCamera��o������NE�,�>�P� �j�|�������ď�I  �v�)��&�8� J�\�n����������ڟ����"�4�[� �vR9˟��������ȯ گ�����"�m�F�X� j�|�����G�Y�I7� ����"�4�F��j� |ώ�ٿ���������� ߳�Y�����Z�l�~� �ߢߴ�[�������G�  �2�D�V�h�z�!߃u nY����������� ��B�T�f�������� ��������Y�"i{�0 BTfx�1��� ��,>P ��Y��i����� ���/,/>/�b/�t/�/�/�/�/cu9 H/�/?!?3?E?W?� h?�?�?F/�?�?�?�?POO/O�j	�u0�? jO|O�O�O�O�Ok?�O �O_�?0_B_T_f_x_ �_1OCO�p�{._�_�_ oo+o=o�Oaoso�o �_�o�o�o�o�o�_ �u���oOas�� �Po���<�'� 9�K�]�o�PEc�� ��͏ߏ����9� K�]�����������ɟ ۟����ϻr�'�9�K� ]�o���(�����ɯ� ����#�5�G�� ;�ޯ������ɿۿ� ���#�5π�Y�k�}� �ϡϳ�Z�����J��� �#�5�G�Y� �}ߏ� ����������������  ��N�`� r�����������<��   $�,� J�\�n����������� ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/��  
��(  }�B�( 	 �/ �/�/�/�/??8?&? H?J?\?�?�?�?�?�?:�*4� �n�O 1OCO��gOyO�O�O�O �O��O�O�O_VO3_ E_W_i_{_�_�O�_�_ �__�_oo/oAoSo �_wo�o�o�_�o�o�o �o`oroOas �o������8 �'�9��]�o����� �����ۏ���F�#� 5�G�Y�k�}�ď֏�� şן�����1�C� U���y��������ӯ ���	��b�?�Q�c� ����������Ͽ�(� :��)�;ς�_�qσ� �ϧϹ� ������H� %�7�I�[�m���ϣ� ����������!�3� E�ߞ�{������� ��������d�A�S� e�������������� *�+r�Oas�������0@  ������� ���)frh:\�tpgl\rob�ots\r200�0ic6_165f.xml�`r �������/����/3/E/W/i/ {/�/�/�/�/�/�/�/ /
?/?A?S?e?w?�? �?�?�?�?�?�??O +O=OOOaOsO�O�O�O �O�O�O�OO_'_9_ K_]_o_�_�_�_�_�_ �_�__�_#o5oGoYo ko}o�o�o�o�o�o�o  o�o1CUgy �������o� �-�?�Q�c�u�����@����Ϗ��K� � 88�?��2��.� P�R�d���������� П���(�R�<�^����r�����ܫ�$T�PGL_OUTP�UT ����/ ���� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ������ˠ2345678901������ ��0�8�����_�q� �ߕߧ߹�Q߽�����%�7���}A�i�{� ����I�[������ �/�A���O�w����� ����W�����+ =����s���� �e�'9K �Y�����a s�/#/5/G/Y/� g/�/�/�/�/�/o/�/ ??1?C?U?�/�/�? �?�?�?�?�?}?�?O -O?OQOcO�?qO�O�O �O�O�OyO֡}�_@)_;_M___q_�]@���_�_� ( 	 ���_�_o�_5o #oYoGoioko}o�o�o �o�o�o�o/U Cyg�����@���	�?��Ƭ� -�G�u���c������� ߏ���`��,�ΏP� b�@��������Οp� ޟ����:�L���p� ��$�������ܯ�X� ��$�Ư�Z�l�J��� ���ƿؿz����� 2�DϮ�0�zό�.ϰ� �Ϡ�����b��.��� R�d�B�tߚ����� �߄�����<�N�� r��&�������� Z�l�&�8���\�n�L� ���������|��� �� FX��|�0 �����d0 � fxV�� ���//�>/P/ �</�/�/:/�/�/�/��/?
2�$TPOFF_LIM [�|�@W���A�2N_SV#0  ��T5:P_MOoN S�74ʌ@�@2�U1ST�RTCHK �S�56_=2VTCOMPATJ8�196�VWVAR rj=�8N4 �?� O�@}21_�DEFPROG �%�:%CON�ROD&O�?_DISPLAY*0�>?B�INST_MSK�  �L {JI�NUSER�?�DL�CK�L�KQUIC�KMEN�O�DSC�REPS��2tpsc�D�A1Ph6Y52GP_KYST�:�59RACE_CF�G �Fr1�4�.0	D
?��XH_NL 2�93��Q�; $B�_�_o o�2oDoVohozj�UIT�EM 2�[ ��%$12345�67890�o�e � =<�o�o�os G !{!@�o ZC�o{�o�� �9K�o/��?� e������#��� G���+���O���ŏ ׏Q�����͟ߟC�� g�y����]������� �����-���Q��u� 5�G���]�ϯ!���� ſ)�տ���q�ϕ� ����3�ݿ�ϯ���%� ��I�[�m���	ߣ�c� u��ρ������3��� W��)��?���ߌ� �ߧ�����c�S�e� w������k����� ���+�=�O���s� EW��c����� �9�o�� n�����#� G�"/}=/�M/s/ �/��///1/�/U/ ?'?9?�/]?�/�/�/ i?�??�?�?Q?�?u? �?PO�?kO�?�O�OO��O)O;O_�TS�R|�_UJ�  �b�UJ �Q`_UI
 �m_�_z_�_8ZUoD1:\�\��Q�R_GRP 1��k� 	 @`@o!koAo/oeoSo�own��`�o�j�a��_�o�o�e?�  '9{#YG}k ����������C�1�g�U�w���	��E��ÏSSCBw 2%[  �!�3�E�W�i�{������\V_CONFIG %]�Q]_��_���OUTPU�T %Y�����S�e�w����� ����ѯ�����+� _A@�S�e�w������� ��ѿ�����+�<� O�a�sυϗϩϻ��� ������'�8�K�]� o߁ߓߥ߷������� ���#�5�F�Y�k�}� ������������� �1�B�U�g�y����� ����������	- >�Qcu���� ���);L _q������ �//%/7/H[/m/ /�/�/�/�/�/�/�/ ?!?3?D/W?i?{?�? �?�?�?�?�?�?OO /OAOݟ�>�O�O�O �O�O�O�O�O_!_3_ E_W_J?{_�_�_�_�_ �_�_�_oo/oAoSo d_wo�o�o�o�o�o�o �o+=Oaro �������� �'�9�K�]�n���� ����ɏۏ����#� 5�G�Y�j�}������� şן�����1�C� U�g�x���������ӯ ���	��-�?�Q�c� t���������Ͽ�� ��)�;�M�_�p��� �ϧϹ��������� %�7�I�[�m�~ϑߣ� �����������!�3��E�W�i�LH�������s���hO�� ����1�C�U�g�y� ��������t�����	 -?Qcu�� ������) ;M_q���� ���//%/7/I/ [/m//�/�/�/�/� �/�/?!?3?E?W?i? {?�?�?�?�?�?�/�? OO/OAOSOeOwO�O �O�O�O�O�?�O__ +_=_O_a_s_�_�_�_ �_�_�O�_oo'o9o Ko]ooo�o�o�o�o�o �o�_�o#5GY k}������o ���1�C�U�g�y����������ӏ���$�TX_SCREE�N 1��;���}��&� 8�J�\�n������ ���ҟ������� ��P�b�t�������!� ίE����(�:�L� ïp�篔�����ʿܿ �e�w�$�6�H�Z�l� ~�������������� � ߗ�D߻�h�zߌ� �߰���9�K���
�� .�@�R���v��ߚ�����������k���$�UALRM_MS�G ?��� ��zJ�\������� ������������/"�SFw+�SEV � �E��)�E�CFG ���  �u@��  A�   B��t
 x�s� 0BTfx�������GRPw 2� 0�v�	 �/+�I_�BBL_NOTE� �
T���l�r��q�� +"DEFPROz5�%9� (%k �/�p�/�/�/�/�/? �/%??6?[?F??j?��?!,INUSER�  o-/�?I_�MENHIST �18��  (� | ��(/S�OFTPART/�GENLINK?�current=�menupage?,153,1�?`O�rO�O�O�)'O9N381,23�O�O�Od	_�O'�O9N71MO�e_w_�_�_*_<ZeditEBCOT_�_�_�oo�A+�_�_ONROD,9#oso�op�o�M&O@_290�_ �o(�_�o�aLO t����B�?�� �	��-�P$�0"A� _�q����������ݏ ���%�7�Ə[�m� �������D�V���� �!�3�E�ԟi�{��� ����ïR������ /�A�Я�w������� ��ѿ`�����+�=� O�:�L��ϗϩϻ��� �����'�9�K�]� �ρߓߥ߷������� |��#�5�G�Y�k��� ����������x�� �1�C�U�g�y���� ������������- ?Qcu`�rϫ� ���);M _q����� �//�7/I/[/m/ /�/ /�/�/�/�/�/ ?�/3?E?W?i?{?�? �?.?�?�?�?�?OO �?AOSOeOwO�O�O� ��O�O�O__+_.O O_a_s_�_�_�_8_J_ �_�_oo'o9o�_]o oo�o�o�o�oFo�o�o �o#5�o�ok} ����T��� �1�C��g�y�����������O��$UI�_PANEDAT�A 1������  	��}/frh�/cgtp/wh�oledev.stmӏ1�C�U�g�R�)pri���]�}��Ɵ؟���� � )"�F�-�j�Q��� ����į���������B�T�;�x�V����   ?  h�F���� ǿٿ����b�3Ϧ� W�i�{ύϟϱ���� �������/�A�(�e� L߉ߛ߂߿ߦ������� ��8���T� Y�k�}������� J�����1�C�U��� y���r����������� 	��-QcJ� n��0�B�� );M�q��� ����/h%// I/0/m//f/�/�/�/ �/�/�/�/!?3??W? ���?�?�?�?�?�? :?OO�AOSOeOwO �O�OO�O�O�O�O�O _ _=_O_6_s_Z_�_ �_�_�_�_�_d?v?4O 9oKo]ooo�o�o�_�o *O�o�o�o#5�o YkR�v��� ����1�C�*�g� N�����o"oӏ��� 	��-���Q��ou��� ������ϟ�H��� )��M�_�F���j��� ����ݯį����7� ����m��������ǿ ����p�!�3�E�W� i�{�⿟φ����ϼ� �����/��S�:�w߀��p߭ߔ���D�V�}����-�?�Q�c�u�)	��ŉ������� ��� ���D�+�h�O� a��������������� @R9v	�`��Z��$UI_PO�STYPE  �`�� 	� ���QUI�CKMEN  ���� RESTORE 1 `��  �i�S`N�m~����� �/%/7/I/[/�/ �/�/�/�/r�/�/�/ j/3?E?W?i?{??�? �?�?�?�?�?�?O/O AOSOeO?rO�O�OO �O�O�O__�O=_O_ a_s_�_(_�_�_�_�_ �_�O�_o"o�_Fooo �o�o�o�oZo�o�o�o #�oGYk}� :o���2��� 1�C��g�y������� ��d����	��-��oSCRE� ?�u1scHWu2h�3h�4h�U5h�6h�7h�8h��USERJ�O�a��TI�j�ksr�є4�є5є6є7є8�ё� NDO_CFG !����Ѩ PDATE ����None� _� ��_INF/O 1"`�]�0%3�x�	�f����� ˯ݯ������7�� [�m�P�������ǿ��J�OFFSET %�ԿσA֏ �*�<�N�{�rτϱ� �Ϻ�Ͼ����A� 8�J�w�n߀ߒ������
����UFR�AME  ʄ��G�RTOL_A�BRT&��>�EN�BG�8�GRP 1�&<Cz  A�����������������:�� U�g��V�MSK  Qj�]�X�N#����]�%�߫��VCC�M�'���RG���*�	��ʄ�ƉD � BH)�p,<2C�)��PN�?�` ��MR��2A0��p���"�р	 ����~XC56# *������N�k�5р�A@<;C� ���ʈ);h�cD��Rр|��Ђ B����6�t/T1/  /U/@/y/d/�/�/�/ �/*/�/	?�/???��c?u?��TCC��1���f�9�ррn��GFS�22w� Й�2345?678901�?�2 ʈ"�6��?!Oс>,1H2�QO_GB@R 8~N:�o=L� ����������O OA�O�O@O_dOvO �O�O�O�_�O�O�__ _�_<_N_`_r_Soeo �_Ro�o�_�_oo&o�8o��4SELEC�F�j�$�VI�RTSYNC� ���6�BqSIONOTMOU-tр���cu��3U���U�(�� _FR:\es\+��A\�o �� wMC�vLOG�   UD1�v�EX�с' ?B@ ����q�DESKTOP-8U37T7F��6��q:�^�σ ��  =	 1�- n6  -#��ʆ�xf,p�#��0=��ʹ����r�xTRAIN���2�1.��
. d��sq4w ( ,1��0��)�;�M�_� q���������˟ݟ����I��crSTAOT 5��@�o�����E:$��ۯ�_�GE��6w�`�. �
��. 2�H�OMIN��7U?��U� �r�a��a�aCG�um�J�MPERR 28w
  ʯE:�� suTs�����߿�� �'�9�O�]ώρϓ�Z_v_�pRE��9t�.��LEX��:wA�1-e�VMPH?ASE  RuC9Cb��OFFLpc�V<vP2�t;4�04�)�8���b@�� x�bb>?s33��Á�1��L��ҕԈ�(|��t�>x��Â�xf�o.���/?P�X� $�2�x���� 0� ���6�+���l� �\�j�|��������� �� �D�V���ZT f���������� . �,BPb� ������/ /(/:/�y/�b/� �/�/L/? ??<? n/c?�/�/�?�?�/�? 6?�?�?�?OX?j?\O �?�OJO�?fO�O�O�O �O0O%_TO_xOm_�O �O�O�_�_�_�__o >_P_EoWo�_xo�_�o�o�o�o��TD_F�ILTEt�?��3 ��Wp��]o$ 6HZl~��� �����)�;��M�_�q������SH�IFTMENU [1@x�<��%�� ��я��0���f� =�O���s�����䟻��͟���P�'�	�LIVE/SNA�PD�vsfli�v�b���I�ON G�U���menu����:������±���A���	0����b�K��5M���U�m`@�����A�p+B8������Ӝ�䝱�����m`� X;ӥ�/�ME��ujY��M���MO���B���z��WAITDINEND�13���OKN�.�'OUT#��Sa�4�wTIM�����GϮ�@���`ϱ����ʞ�2�RELEAcSE����TM������_ACT�x��Ȫ�2�_DATOA C�ի�%i�x�ߪ���RDIS�~b��$XVR2��D��$ZABC_GRP 1E8��n`,@h2��ǽZIP1�FD� cCo�������x�MPCF_OG 1G8�n`0<o� ���=�H8����t�� 	�w�  8R�����e�����?�k������5���
\��  �a �����7�����I��z��_YLIND�aJ��� �f ,(  *s�K�p���� �// +.mN/�r/Y/k/�/ ��/�/�/3/?�/�/ J?1?n?U?�/�?�?v��C�2K8��� � �O`o�7O~[Olh�?�Og��AA�A�SPHERE 2LS�?�OX?�O_ _>_�?�Ot_�_?�_ I_/_�_�_o�_]_:o Lo�_�_�o�_�o�o�o��o#o $7�ZZ� �k�