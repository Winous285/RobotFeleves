��   u��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����UI_CONF�IG_T  �� A$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]2�ODE�
3CWFOCA �4C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"��%�!BA�!j ?Ɵ"BG�%�!jIN=SR$IO}7�PM�X_PKT��"IHELP� M{ER�BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�; } &USTOM0� t $} R?T_SPID�,D�C4D*PAG� ?�^DEVICE�PISCREuEF���IGN�@$FLAG�@C�1 � h 	$PWD_ACCES� E �8��C�!~�%)$LABE� O$Tz j�@��3�B�	&U�SRVI 1  < `�B*�B�n�APRI�m� �t1RPTRIP�"m��$$CLA�@ ����sQ��R2��RhP\ SI�qW�  �
�QIRTs1q_�P�'2 L3hL3�!pR	 ,���?����Q�P�R�T�Q���S���P�  o��
 ��zQQoco uo�o�o�o�o Mo�o �o*<�o`r ����I��� �&�8�J��n����� ����ȏW�����"� 4�F�Տj�|������� ğ֟e�����0�B� T��x���������ү a�����,�>�P�b���PTPTX���򨅿���P �sm���$/so�ftpart/g�enlink?h�elp=/md/�tpmenu.dgd����"�4��X� j�|ώϠϲ�A����� ����0߿�A�f�x� �ߜ߮���O�������,�>����zQ�'`V�	bbS� ($ �ߕ�����������zQ�Q�c����I��k
m�d����
a����  ���	����@�d�n���	f�P#` � �V������SB �1�XR �\ }%`;REG VED��� wholem�od.htm4	s�inglEdo�ub\tri�ptbrows�@�!���� /AS|�|/Adev.sJ�l�o�1�	t ���w�G/Y/k/�5/�/�/�/�/�/ ?� �P?*?<?N?`? r?�?�?�?�?�6�@? �?�?�? O2ODOE	 �/�/wO�O�O�O�O�O �O�O__+_=_O_a_ s_�_�_�_�_��_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -??z��� ����
��O@� R�!�3�����QOcOI �ݏ��*�%�7�I� r�m��������ǟٟ �����_/�)�W�i� {�������ïկ��� ��/�A�S�e�w��� ��iֿ�����0� B�T�f�x�s��Ϯ�}� �����ϭ�����>�9� K�]߆߁ߓߥ����� ������#�5�^�Y� k�9����������� ����1�C�U�g�y� ��������������ſ 2DVhz��� �����
��@ R	������ ���/*/%/7/I/ r/m//�/�/�/�/�� �/�/?!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSO!�O�O �O�O�O�O�O__0_ +T_f_5_G_�_�_�Z��$UI_TOP�MENU 1��P�QR �
d�QfA)*defaultqO�ZM*leve�l0 *\K	 o� So�_Qocb�tpio[23]��(tpst[1��heo�ouo3oEo�-
�h58E01.g�if�(	mencu5&ypHq13&z�Gr%zEt4M{4�a��������� eB�C�U�g�y�����~,�prim=Hq�page,1422,1��ݏ��� %�0�I�[�m�������2���class,5������)�4���130�f�x�Њ�����5���53�ʏ���� �2�5���8ٯm�������� 4�ٿ����!�3�^I�P�Q�_k�m]��a0[ϕ�o�fty�m�o��amf[0�o��	>��c[164�g.Ճ59�h�a���tC	8$|Gr2uK}��az mWw%{�ߩsK�]�6� H�Z�l�~�ɿ�����`�����𢡊��80$�?�Q�c�u�����̐2 ����������	��ʟ ?Qcu�(T��������Ѥ1�.�N`r����~��ainedic�����//��c�onfig=si�ngle&��wintpĀ /`/r/�/ �/]J�QV¤/�/e�/ �o�o??1?D?U?g? y?�?�/�?�?�?�?�? 	OO-O?O�aO�O�O �O�O�O�O��__*_ <_N_`_�O�_�_�_�_ �_�_m_�_o&o8oJo \ono�_�o�o�o�o�o �o{o"4FXj �o|������ ��0�B�T�f�x���������ҏ���MN S�,�wω¯����w����s��<����ϡ�u0�͔�V�|�F7��7�����԰�Οp��ߔ�6��u7��� ����`�/�A��227� ��������˿Z�l���@��,�>�P�/!$13�ϛϭϿ��ϐ� ����+�=�O���s� �ߗߩ߻�����"�߀�'�9�K�]�����6 d��������,$۬74r��/�A�S�e��,����%	TPTX[209�����24����������18�������
����0P2���1_��E�tv�����Q�u10�1=�ïqC�:4$treevi�ewA#�3�&d�ual=oU81,26,4��� �n����	//-/ �Q/c/u/�/�/�/ֺ	;@b�3`r�? )?;?F/_?q?�?�?�?��?�/�/\2�/t2@��O1OCO�?��1�/`E���O�O�O�6XO��edit�zO�O _._@_׹?���OC L_�_�_�_~��_�_G� o}o�CoUogoyo �o�o�o�o/o�o�o	 -?Qduӥ� ������I?2� D�V�h�z������ ԏ���
����@�R� d�v�����)���П� ������<�N�`�r� ����%���̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� �_�_X�o|��o��� �����������ߋ� )�S�e�x߉ߛ߭߿� �ߓ��,�>�P�b� t￿���������� ���(�:�L�^�p��� ������������ �� $6HZl~� ������ 2 DVhz��� ���
/�./@/R/ d/v/�/7�IϾ/m��/ I���??)?;?M?`? q?�?�/�?�?�?�?�? OO%O7O��nO�O�O �O�O�O�O%/�O_"_ 4_F_X_�O|_�_�_�_ �_�_e_�_oo0oBo Tofo�_�o�o�o�o�o �oso,>Pb �o������� ��(�:�L�^�p�� ������ʏ܏/�/ $��/H��?MOk�}��� ����ş؟�W���� 1�C�U�h�y�����_O ԯ���
��.�y�@� d�v���������M�� ����*�<�˿`�r� �ϖϨϺ�I������ �&�8�J���n߀ߒ� �߶���W������"� 4�F���X�|���� ����e�����0�B��T���*def�aulta�2�*?level8��������{� t?pst[1]���ytpio[#23��u�������	menu_7.gif�
�13�	�5�
��
�4�u6�
ʯ? Qcu����� ��//�;/M/_/�q/�/�/�/6"pr�im=�page,74,1�/�/�/�??+?6"�&cl?ass,130?f?@x?�?�?�?=?O25�?@�?�?O O2O5#D< �?lO~O�O�O�O�/�"18�/�O__'_9_DON26@_u_�_�_�_��_��$UI_U�SERVIEW �1��R 
���_>��_
o�m(oQoco uo�o�o<o�o�o�o�o �o);M_qo ~������ %��I�[�m������ F�Ǐُ������ .�@���{�������ß f������/�ҟS� e�w�����F�P���̯ >���+�=�O�a�� ��������Ϳp��� �'�9��F�X�j�ܿ �Ϸ������ϐ��#� 5�G�Y�k�ߏߡ߳� ���߂������z�C� U�g�y��.������ ������-�?�Q�c� ������������� )��M_q� �8������  2�m�� �X���/!/3/ �W/i/{/�/�/J�/ �/�/B/??/?A?S? �/w?�?�?�?�?b?�? �?OO+O�/�?JO\O �?�O�O�O�O�O�O�O _'_9_K_]_ _�_�_ �_�_�_lX