��   ��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A 	  ����DRYRUN_�T   � }$'ENB 4 �NUM_PORT�A ESU@$STATE P _TCOL_��PM�PMCmGRP_�MASKZE� O�TIONNLOG�_INFONiA�VcFLTR_E�MPTYd $P�ROD__ L �E�STOP_DSB�LAPOW_REwCOVAOPR��SAW_� G %$INIT	�RESUME_T�YPEN &J_�  4 $�($FST_ID1X�P_ICI0 �MIX_BG-yA
_NAMc �MODc_US�d�IFY_TI��.yMKR-�  $LIN�c   �_S�IZ�w� k. �, $USE_FL4 ��&i*SIMA�Q�#QB6'SCAN��AXS+INS*I���_COUNrR�O��_!_TMR�_VA�g� h>�i) �'` ��R��!�+WAR��$}H�!{#N�PCH��$$�CLASS  O���01��5��=5%0VERS�.7�  �=
A1IRTU� .?�@0'/ l55�������Y0�6!m071�5��%71�?����?
O��}5I2�;�GOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_��%FW�?N8�0 @���_J�[m0�]�o �{ 2�; 4%t_$o���1�1o Wo6o{o�olo�o�o�o��o��8�o��G"q 
O��= ">���" wry�S�P��=�9Y0���t�1�tX�1l1Y0�> �&�8�J�\�n����� ����ȏڏ����6�1 ��1 �2�D�V�h�z� ������ԟ���
��44�6�S!2�9 �[�m�� ������ǯٯ���� !�3� �M�f�x����� ����ҿ�����,� >�I�b�tφϘϪϼ� ��������(�:�L� W�p߂ߔߦ߸����� �� ��$�6�H�S�e� ~������������ � �2�D�V�a�z��� ������������
 .@Rdo���� ����*< N`k}���� ��//&/8/J/\/ n/�V