��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�   � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d PPINFwOEQ/ ��L A �!�%/� H� �&�)EQUIP 2� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CESS0s!_81s!J3�> �! � �$SOFT�T_�IDk2TOTAL7_EQs $�0�0�NO�2U SPI_OINDE]�5Xk2SCREEN_(4�_2SIGE0�_?q;�0PK_FI�� 	$THK�YGPANE�4 �� DUMMY1"dDDd!OE4LA!�R�!R�	 � �$TIT�!$I��N �Dd�Dd ��Dc@�D5�F6�F7*�F8�F9�G0�G�G@JA�E�GbA�E�G1�G( �F�G1�G2�B!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HO30IO�0� }%�SMACRO�ROREPR�X� D+��0��R{�T UT�OBACKU��0 �)DE7VIC�CTI*0�A� �0�#�`B�S�$INTERVA�LO#ISP_UN9I�O`_DO>f7�uiFR_F�0AI�N�1���1c�C�_WAkda�jOF�F_O0N�DEL��hL� ?aA�a1bc?9a�`C?��P��1E��#sATB��d��MO� �cE' D [M�c���^qREV�BI�Lrw!XI� QrR�  � OD��P�q$NO�^PM�Wp�t�r/ "�w� �u�q�r�0�D`S p �E RD_E�pCq�$FSSBn&$CHKBD_SE^e�AG G�"$SLOT_��2=�� 	V�d�%��3 a�_EDIm  O � �"��PyS�`(4%$EP�1��1$OP�0�2��a�p_OK�UST1P_C� ��d���U �PLACI4!��Q�4�( raCOM9M� ,0$D�����0�`��EOWBn�IG�ALLOW� �(K�"(2�0VAARa��@�2ao�L�0;OUy� ,Kva�y��PS�`�0M_Ox]����CF�t7 X� GRP0�z�M=qNFLI�<ܓ�0UIRE��$�g"� SWITCH^ړAX_N�PSs"�CF_�G� }�� WARNM�`0#!�!�qPLI�I�wNST� COR-�0bFLTRC�T�RAT�PTE�� $ACC1a�N ��>r$ORI�o"v��RT�P_SFg� CHG�0I���rTא�1�I��T�I1��� x� i#�Q��HDERBJ; C,�2'�U3'�4'�5'�6'��7'�8'�9{5CO`T <F П���x�#92��LLECy�}"MULTI�b��"N��1�!���0T_�}R  4F S�TY�"�R`�=l�)�2`�����`T |� �&$c�Z`�pb���P�MO�0�TT�OӰ�Ew�EXT�����ÁB���"2�� ��[0�]�}R���b�}� D"}����Q���$Q�kcG���^Ȉ�1��ÂM���P��� ŋ� L@�  ���P��`A��$JOBn�/�i�G��TRIG�  d �p�߻���³�7��4�����_M�b�! t�pF� CNG AiBA� ���� M���!���p� �q�ᄅ0��P[`��i�*�"6���0tB񉠚�"J��_Rz�gC��J��$�?�Jk�D�%C_�;������0Ф}R�t#� ��ȩ���G���0NHwANC̳$LGa��B^a��� �D��!A�`��gzRɡ�!`��p�DB�fRA�AZ�0�KELT�Ė��PF+CT&��F�0�P&��SM��cI��1 �% ��% ��R��a���� S��&����M 00{o e#HK
~�A^S��������I_T$�"6SW��CSXC)�?!%���p)3��T�$�@��PANN&�AI�MG_HEIGH�Cr�WIDI AV�T�0��H F_A�SPװ��`EXP��1���CUSTJ�U��&��|E\�!%�C1NV _�`�a���' \%1y�`O�R�c,"�0gsk��PO,��LBSYI�G��a R%�`좔Pspm��0k��DBPXWORK���(��$SKP�_�`ma�"<qTR>p ) ���P`���� �0�DJ!d/�_CN��R�#� �'�PL�S�Q�d�s�DKA7WAw'�^A0�@NFZpfBDBU��*�"!PRS�7�
pЖQ����+ [pvr�$1�$ZϢ�Li9,v?�3ʠ��)-�?�4C��.�?�4�ENEy��� /��?�3J0RE`��20�H��CuR+$L,C,$i3
�? =KgINE@�K!_D�I�RO�`����ȳ`qvC��h �FPAÃ�3uR�PRN�B�MeR��U!�u�CR[@�EWM �SIGN��A� .q�E�Q�-$P��.$�Pp 2�/ P7�PT2�PDu`L����VDBAR@�GO_AW���Jp � ��DCS�pZ�CY_' 1���@1<�Q�?fIG2�Z2>fN�>�����
�qS&c}P2� P $��RB�?�e�P=hPwg�QB�Yl�`gT+1�THNDG�23��KS�SqE|�Q��SBL㠸�cc�T�qSL��4 HpZ ���VTgOFB�l�FEfA��ǿb�TqSW5�bDqOC���MCS�f��`Z$r�b H� W�0��T�"sQSLAVv�16�rINP���f��LyqQP�7� $,�S���=���v��uFI���r줭sc�!��!W�1ԭrNTV'��rV�	��uSKIvTE��@W���:�J_� _�00�SAF�E�A�_SV��EOXCLU��B �P%DJ L1�k�Y�d�Ɯ�rI_V� !P�PLY 0b���DE�~w��_ML2�B ?$VRFY_�#��Mk�IOU��憻 �0���:�O�P��LS�@jb;�3572��S	r�� Px%X�{P�8hs� �� 8 @� �TA� qঠ ��c_SGN��9 6����@�A�����i�Pt!��s"��~UN��0jdՔ�U���B  �@� ��� ���K�t�W I�2: @�`1Fؒ���OT�@@Ð:41(�774C2�M`NI�2;�R����r��A�q��DAY1#LOAD�T/4~�;3�0� �EF�XIJ�b< @%1O�|�3� _RTRQ��G= D�`@��Q@  �EjP"�㥂��<�B�� 	�@��GAMP��]>��a�����a�8Sq�DUt�@q���"CAB���?A��0NSs���IDI�WRK�^�� �V�WV_]���> ��DI��q�@�� /.�L_SE2�T���/�Z`��0��#�E_��u�v�j��SWJ�j� 𐲰��	���=c�O�H�z�PPJ�v�I	R!��B� ��w�d�p�B"����BASh���� X ���V����?�C��Q��RQDWf��MS���AX}�<8�u�LIFE� �7�A1C�NJ���S��DH���Cs�>��C`QN"�U��3OV� _�HE����'SUP�hbC�� _�Ԥ���_����[Q
��Z��W���ו�Tb��XZ$ `1��+Y2F�CM@T��t@�N�p��!��9gA `�P.�HE��SIZy֥�u��B�N�pUFFI����p� �Q/40�<26�71#�!MSW9B� 8�KEYIMAG�CTM@A���A�Jr��!OC�VIET���C �C�V L�t���s?�� 	�!� :D�6"pST�!x�0��� 0��Ѡ��0���EMAIL���@�����c`_FAUL��E8H�CCOU�p}$�T@��F< �$���eS]���ITvBUF��q���T�  ���BdC�t����#��SAV b$)�e�A� }����Pi�e@U�b`_0 H���	OT{BH��lcPր(0�
{��A�X1#�� @��_9GJ�f1YN_�� EGj�D�U/0e��UM����T8�F���ِ�A!H�0(@u���C_r@�@AK�D����=pR�8���uDSP �uPC�IMb��J���U��ЁEƀF��IP�su��D`��TH0�c��T�uA�HSDI�AGBSC�ts��0Vzp�*} �$�#��NV�W�G�#�$0� F�J�/d�j�ASqC��U�MER��>uFBCMP��t�ETH�!AI��FU��DU �a�@;⠂�CD�O � ���R�_NOAUTg` J��Pp2��n4VĥPSm5C`}5	CI�.2qk3� =_KH *}1Lp ��Q��&�I���4 #Q�6s��6ѡ�60��6T���67�98�99�:�J��8�:1J1J1�J1+J18J1EJ1*RJ1_J2mJ2�;JU2J2J2+J28JU2EJ2RJ2_J3mJ%3�:3KJ3J/�TG8J3EJ3RJ3_J94mB|�EXT�>aLC`��F�fF�5pQ9g�5��FDR�/MT��VC��pC�wa}"C�REM,�9FAj�OVM��e�A�iTROV�iD�Tm �jMX�lINp�i���j�IND�`�!�
xp /$D�G���`opS�9�D��`RIV)0Qbj�oGEAR�IO0�	K�bu�Nj�x�.�����p�qj�Z_MCaM>�C�d`��UR)2�N ,{1��?� ��
 ?�pI�?�qE���q��T�0lbO����P�� �RIT5��UP?2_ P Ѡ#TD= ��C����qP��J��0.�BAC;QC T��$9 O�)��OG��%E��3e&0IFI��e0�0��梅PT��1FMR}2ieR vbY�vbLIq��{g�����f��Ŗb_mAN~F�_F�I4+��M;v`r}DGCL�F��DGDY��L�D�q>t5[�5S��$ہk�SY�M�� T�FS� l�T� P�)���
�/�$EX_)�@�)�1P�� ��*�3b�5b�s�G�!ieU � p�&2SWKO��DE�BUG�S��0�GRtY�zU�#BKU� �O1�@ O�P�O8��Π0��ΠM�S]�OO��SM�]�Eq��pQ`_?E V $�o��TERM2�W;�� �ORIĀ6�X~;� �SM_���$7�Y;�`��TAry�Z;����UPB�[� -��Qb�V$G���W$SEyGźאELTO���$USE0NFI����p���`�>��X$UFR����`q0豈�D5h�OT1�ƴ TA_ �C�NSTd�PATT!��Y�OPTHJ!B0En�8�K0�ART� ��p������REL��&SHFTF"�_�.��_SH��M�!B0"x� ��n���Z����OVR
#&SHIԾ���U�2 �AY#LO$ 5I1�p_�d���d�ERV�0 *�} ��b?�d��Q0����A��RC
���ASYMh���WJ�apE�����f�2�U��d�5����D5��P#Gи!	�OeRd�M��GR!���\��΢�^��8���k�] �E�]��TOC���q��OP��N z�3�&1���aO�a> R%E��R�#&O0��`�e��R]�����|����e$PWRSp3IM��[�R_����VISy�r���UD��t�� ^>��$H����_ADDR9fH$�Ga�z��s�i1R� =_ H8�S� ��S��C0��C��CSE�a�baHSO0��` $���_D`����PR�vt�TT� UTH��a ({0OBJE�1u���$9fLE�P�-=b � �*g!AB_qT���Sk�#DBG�LV5#KRL"�H�IT�BG0LO:���TEM4$�0�b������SS�p�4�JQUERY_FLA��f WYA���ec��� PU�"B�IO0��4G���H��HB �IO�LN~�d/0i�C^��$SL�� oPUT_�$���Pwp�rSLA�� e/2�����ӡ�ҽ1IO F�_AS�f��$L��U���#�04�#0����,�HYOgN!�'#�UOP�g ` l!9f�b>$�`E&�!��P����'�!E&��"�&�P_ME�MBk0T h �X IPz�v��"_ #0v����0��Oc6��1w�DSP�' $FOCUSBGv���0UJhfi � 860S��JOG�W2�DIS�J7��O^��$J8�97���I6!�2�77_LA�BQ����0�8�1AP�HI�pQ�3�7D�+�J7JRA4`P�_�KEYp ��KILMON�j&`$XR =0c?WATCH_ �D�L��U1EL� �y`LB�k GpG�VP�-ffBCTR��fB5vbaLG|�l ���+h�"��LG_SIZ{Y��E
��F
 �FFD�HI�H�H��F �HM��F�@���C5V
� 5V
 5V�@5VM�5W�`AS)@S����@Nv1
��mx � ��R���4a�PÀU�Qk�LܲS�RDAU�UEA` I���R�PGH���؁ BOO~�ng� C-"2�ITGc�d��)&REC-jSgCRN)&DI(#S��RG����cl@�!#��b�!Sa�"Wkd!�T!#JG=M�gMNCH"�FN�2�fK�gPR�G�iUF�h	��hF�WD�hHL/ySTP�jV�hĀ�h`�h�RSgyH!�{&C��Es��!#���g�yU t�g�¬f|@6#�bG�i4�PO�JzZebEsM�w82�iEX'�TUI�eIP�c w��c���c���`�a�����s��Jg��KaNO�{�ANA"貇�V3AI�0zCL����?DCS_HI���������O����SI�)��S'��hIGN �@��C�aT����7DEV�wLL�єQ�6@BU𠔠oa@��T��$�GEM�'9nDcѢ��p�a@ЅC�!��O+S1��2��3��d9_����q �T0v�-�絡.e�IDX����-fL�b�STm R�PY0����� p$E��C ���  ����� ��r L*</��Q(06����6�EN 6��ՕKc_ s �Y��P$ dKaD� �{MC�Rt �T0�CLDPm ��TRQLI`��e0x�f��FL>1��_����DUA��LD������ORGe0�r���WX������Y���V�O�u � 	���uu���%Si�Tx��00�ް�S�[�RCLMC�i����{�m[�ՐM9I��O�v d�Q6��RQ�00�DSTB��Y� ��{a���AX��@�� �EXGCES�����M�
��wA0�¹�+�j��x(��_A�ʠ� l����V�K|�y� \*�2��$MB�LIE��REQGUIR����O��ODEBU��L�M{�zW�.!��B�ӊi���N,03Ѩ�{0�R�RkHV�DCE��T�IN3 `!�TRSMw0p�S�N�����s<�wPST�  |h�7LOC9�RI� 9�EX��A��:������ODAQo%}��1$@�Q΂MF�A �_���p�C��P���SUP�ՐFX���IGG�"~ �0��MQ���v�5@� %����m ��m x����6#DATA�����E� 1�NP" Nn�� t�MDIF)?�!���H���1!� �1"ANSW�a!ܑS�!�D�)��H3Q�$�[ ?�CU�@V_ �>0���LO�P$�H=ұ���L2��t����RR2I5��  ��QA�X� d$CALII��NUG�2g�RINp<$R�SW0��K�A�BC�D_J2SqE����_J3v
p1SP�@6 ��	Pp�3��\�����J���P�O村IM��[�CSKAP��$�P�$J�Q[�Q,6%%6%,'���_AZW��h!ELx�����OCMP�����1X0RT�Q�#�c1�c@�Y�1��(t�0�*Z�$SMG�p�����ERJ�ԑIN� ACߒ�@�5�b��1�_B��542d���14X҆f>9DI~!��DH �t30���$Vlo�Y�$�a$�  ��A�<�.A�����H �$BE�Ly lH�ACCE�L?��8���0IR�C_R��0�AT<w�c�$PS �k�L  �0F��0Gx�Q�FPATH�9�WG�3WG3&B��#�_@�2�@�AV���C;@��0_MG|a$D�D�A@[b$FW�(����3�E�3�2�HD}E�KPPABN.GROTSPEE�B���_x�,!��DEF�g��1&@$USE)_��Pz�C ����YP�0V� �YN���A{`uV�8uQM�OU�ANG�2�@O9LGC�TINC~����B�D���W���ENCS����A�2��@INk�I&Be���Z�, VE�P'b2�3_UI!<�9cLOWL3��pc x��UYfD�p��Y�� ��Ury�C$0 fMOS`�Ɛ�MO����V�PE�RCH  vcOV�$ �g9��c��\bYĀ���'�"_Ue@0��A&BuL������!epc�\jWvrfTRK�%h�AY�shчq&B��u�s���&l��Rx�MOM|���h�ﰞ �Ą�C�sYC���0D�U��BS_BCKLSH_C&B��P �f�`}S�7��RB��Q.%CLAL��b?�8�pX�t�CHKx�H��S�PRTY�����e�����_~��d_�UMl�ĉCу�ASsCLބ PLMT��_L�#��H�E ������E�H�`-��Q#p_��hPC�aB�hH��ЯEǅCw���XT�0�GCN_b(N�þ���SF�1�iV_RG�e�!��&B����CATΎSH ~�(�D�V��f�0'A�	� �@PA΄�R_Pͅ�s_y�뀎v`�`x��s����JG5��6Ф�G`OG���rTORQUQP��c�y��@�Ңb�q�@�_W �u�t�!�14��33��3�3�I;�II�I�3F��&������@VC"�00���©�1��2�8ÿ�¶�JRK�����綒 DBL_SMt�QO�Mm�_DL�1O�GRV:�3ĝ33��3�H_��Z@a��COSn˛ n�LN ���˲��ĝ0��� �� e��ʽ̃��Z���f��MY���z�TH|��.�THET0beNK23�3Xҗ3��[CB]�CB�3C��AS���e��ѝ3���]�SB�3��h�GT	S@! QC���'y�x�'����$DU�� ;w	��Q�����q9Q����$NE$T�!I�����)I7${0LсAP�y��`�k�k�LCPHn�W�1eW�S�� �������W���������{0V��V��0��UV��V��V��V��UV��V�V�H��@����7�����H��UH��H��H�H��O��O��OF	��O���O��O��O��O*��O�O��FW�}���	�����SPBA�LANCE�{�LmE��H_P�SP1��1��1��PFULC5\D\��:{1��!UTO_���ĥT1T2��22N���2, ����q^P<�-B#�qTHpO~ |�1$�INSEG�2�{aREV�{`aD3IFquC91�('o21�dpOB!d�=���w2��7P���LC�HWARR�2AB����u$MECH`��ДQ�!��AX�q�PB��&r�~2�� �
�"��1eROBƬ`CR&B�%��J?�MSK_�4_� P �_OPAR�1�2(47Qst1��,`*R(0)cB�(0|!I�N!�MTCO�M_C���0� � �@0 �A$N'OREc�2�l ~2o� 4�GR��%FLA!$XYZ_DA��LP;@/DEBU�2 �0lR֫0� ($mQCODS� �2�r� ��p$BUFI�NDX*P �2M{OR3� H%0 �p�0��:@�p�QB�"��1��NF�TMA9Q#C�rG.B�� � $SIMUL���0�As�A�sOBJE3�FA�DJUS�H�@AY�_I��xD�GOU�TΠ�4�p�P_FI�Q=8AT#�Y,` W�1P +�PQ+ 9�:uDjPFRI �PUMT0�RO�
`E+�>Sp�OPWO��0��,@SYSByUi� @$SOP�Q�By��ZU�[+ PR�UNn2�UPA;0D�V�"�Q�`_�@F��P�P!AB�!H��@IMKAGS�%0?�P!3IMQAdIN$��R~cRGOVRDEQ�R�@�QP�Pc�� �L_��feÂސR�Bߐ<pX�MC_SED'@�  H�Ni �M�bG��MY19�F�#@EaSL30�� x $OVS�L�SDIsPDEAXǓ�f֓Hq�bV+��eN�a
��Pp�cw�x�bw�
�d_SE9T�0� @�CrL�%9�RI�A3�
Vv!_��bw{qnq#@-!\�@� �4BT� �àATUS�$�TRCA�@PB�sB�TM�w�qI�Q�d4pF��s�`0� D%0!E�P�b�rr�E1"�qpQpd��qEXE�p@���a�"��tKs�Rp�&0�pUP�01�$Q `XNN�w���d����y �PG|5�� $SUB�q�%xq�q|sJMP�WAI$�Ps��L�O ��1
 �E$R�CVFAIL_C@1�PÁR%P�0�#����Ȕ� �
�R_P=L|sDBTBá��ΧPBWD��0UM��IG�Q `�,�GTNL ��b�ReQ��2���qP��@E�Ǔ��֒��DEFS}P� � L%0ĺ ��_���CƓUN!I�S�wĐe�R)���+�_L
 P�q�#@PH_PK�5�~�2RETRIE|s̛2�R���FI~�2� � $��@� 2��0DB�GLV�LOGSCIZ�C� ���U��2|�D?�g�_T:��!eM�@C
 #EM���R��y0�8CHEC�KS�B�Po01�B�0.�0R!LbNMGKET��@�3砹PV�1� h�`A�Rp� �1)P�2>�S��@OR|sFORM3AT�L�CO�`q�d���$Z��UX�P�!r:�LIG�1� w ˣSWIm ��a#@��,�G�AL?_ � $`@R��B�a��CS2D�Q�$E1��J3�DƸ� T�`PD�CK�`�!LbCO_J3����T1׿6� �˰C_Q�`� � ��PA�Y��S2u�_1|�2|�ȰJ3�ИˈŬƼ��tQTIA4��5:��6S2MOMK@�à��������y0B׀A�D��������PU��NR��C���C����?q��4�` I$PIN�u�41�ž� ��:q�R~ȇ��ٯ� �:�h��a�֬��ց��1�'1R\uSPEED G��0�؅�� 7浔؅�%P7�m�F�p�U��؅SAM �=G��7��؅MOV	B� e0�� ��c2 ��v��浐�� ���c2@nPsR����İ$QH���IN8�İ��?�[��6�؂A���X����G�AMM�q�4$GGET1R@�SDe�zmB
�LIBR[��y�I�7$HI�0_�5a@c2E`@#A@ 1LW^U�@	�1a¬&o�ʱC�=�n S`�p �I_��pPmDòv� ñ'����mD��	ȳ� �$�� �1��0IzpR� D`T#|"c���~ LE^1�41�qwa�?�|�M�SWFL�MȰSCRk�7�0��Ѻpv���Z 0�P�@�9@���2�cS_SAVE_Dkd%]�NOe�C�q^�f�  ��uϟ�}ɕQ��}��Ѐ}*m+��9��ժ(��D �@���������b3 1�RA�Mam�7
5�#���^���Mtա 7� �YL��
A
'�VAS	BtRna`7 GP�B
Bl3
A%`�$GSB1W? �2�2c�Ȭ3oBB1M&@�;CL �8���G�b�1v���9M!Lr� �N�X0�d$W @�ej@b �� @=�BD�BK�B �-�> �P����ycJİX �OL�ñZ�E����uԣ ��OM�R/d/v/�/ �/��A�jM`��e�_��� |��H  ��jV��yV��yP�ʗW�V��E�����NR������NTP=���PMpQU�� �� 8TpQCOU�,�QTHQ�HO�Y2`HYSa�ES���aUE `"#�O.���   �P�0��rUN�p�3��O$�J0� P�p^e��x����OGRA�q�k22�O�d^eITxm�aB`INFOI1����k�ak2��O�I�b� (!SLEQ(��a��`�foayS� ��� 4Tp�ENABLBbpPTION|s����Yw���1sGCF��O�c$J�ñfb����R�x!�]ot vq_sEDŀJ0� �N�R�@K�᪃ES sNU�w�xAUT,!�uCOPY�����v�8 MN����PRUT�� �Nv�pOU��$Gcb|n���RGADJI1ͮ2�X_B0ݒ$P ����@��W��P��`���@㊀��EX�cYCLB����NS6u9�N0�LGO�A��NYQ_FREQ�Z�W���+�p�\cL�Am"����Ì�uCcRE  c� IF�Ѷ�cNA��%i�_}GmSTATUQP<mMAIL�� 1���yd����!��EwLEM�� �7 >DxFEASIGq2 ��v��q!�er$�  I�`�"��ae�L|I�ABUq�E�`rD�V֑a�BAS���b� [�Ub�r % �$y���RMS_TRC�ñj���Ca����ϑ��,r���C��YP	 � 2� g�DU�����Ԣ��0-�1��1���qD�OU�ceNrs��P�R30;p�rGRIyD�aUsBARS(�sTYHs��OTO�RI1��P`_��!ƀ䬲l�O�@7t� �s �`�@POR�c�ճ��ֲSRV��),���DI. T����!��+��+�4)�5*)�6)�7)�8��a�F��:q�M`$VALU|�%�ޡ��>7t�� Cu'!ğa���� (gpAN�#��R�p0� 1T�OTAL��[��P�W�It�&�REG#EN$�9��SX��sc00��Q���PTR��Z�$�_S ��9дsV ���t���rb�E��x��a�"^b�p��V_Hƕ�DA�C����S_�Y4!�B<�S�AR��@2� f�IG�_SEc���˕_�b`��C_����w���?r��%�b�H�SLG#�I1��p"=����4��S�2̔DE��U!Tf.p��TE|�@���� !a�����Jv�,"��IL�_MK��z�н@T�Q�P�a����2V�F�CT�P���^�M�u�V1t�V1��2���2��3��3��4��4����С����1�"IN	VIAB@N�; �!B2>U2J3>3J4>�4JI05���"���{p�MC_F`3 � L!!�r��M= I��M� �[PR�� KE�EP_HNADD"�!f�C�A��A!����"O�Q  I����"��?�"REM9!�ϲ�^uzU��e!HPWD  _SBMSKG�a�	!B2B�
#COLLAB�!��2��h���o��`IT�p�A`��D� ,p�FLI@��$SY�N� ;,M�@C>��~%�UP_DLYI1=�MbDELAm �ژ�Y�PAD�A��`QSKIPE5�� ��``On@NT�1� P_``�b�' �`�B]0�'���)3��) ��)O��*\��*i��*�v��*���*9�JS2R‎��?sX��T%�|1�{2ܐ�p|1�a��`RDC!FW� ��pR�sR�PM�'R^��:b�2��RGE�p2��3d�F�LG�Q�J�t�SP9C�c�UM_|0��_2TH2NP�F@~o0 1� �0�EF�p11��� �l[P�E-Ds#AT Wo�[�w�B�`�d�A �p3�BfcAHnP�B��_D2gB�mOO�OP�O�O�O�G3gB��O@�O_ _2_D_�G4gB�g_y_�_�_�_�_�G5gB��_�_oo,o�>o X_D6gBŀaoso�o�o�o�o�G7gB��o�o&8
�G8gB�[m�H���ES����\@ǡ`CN�@K_@w-E��^� @o�L�m�IO�ፉI���Г!R�@WE!� W�: �1���0�� �5%Ȃ$D�SB;���֒ �h C�L@���1S232Ns�� ��0�u.���ICEU{���P�EV@��PARIT��њ�OPB ��F7LOW�TR2��X�]���CUN�M��UXTA���IN?TERFAC3�f�U��	�CH�� t� � ˠE�fA$����OM���A�0נI���/�IA�TN���T�p� ��ߓ��EFA� p�"!�Ґ�� u!$��� O�� &*��� �����  ?2� �S�0�`?�	� �$3@}%!:B�Ŏ��_���wDSP��JOG���V�h�_P�!s�ON�q0%�0���K��_�MIR���w�MT7��AP)�w�>@"����;AS������;AP=G7�BRKH����G �µ! ^���i����P��Ҏ���BSO�C��wN���16��SVGDE_O�P%�FSPD_OKVR�u �Dв&ӣOR޷�pN��߶�F_�����OV��S!F�<��
�F0�����UFRAF�TO�d�LCHk"%�OVϴ ��W[ ����8�Ң�͠;�  �@ BTIN����/$OFS��CK��WD���������r����TR��T�_�FD� �MB_C �B��B����(�.Ѻ�SVe���Ȅ�}#�G)�<�AM���B_��jթ�_�M@�~��ቂ��T$SCA����De����HBK�����IO���թ���PPA ��������Տթ���?DVC_DB��?� ���A��,�X� b���X�3`���3�0��Ć�ϱU󳠈�CAB�0��ˠ��c� ��Ow�UX��SUB'CPU�ˠS�0�0 �R����!�A�R�ł~�!$HW_Cg@ A��!��F��!�p� N� �$U r�l�>e�ATTRI��y��ˠCYC����CA���FLT ���������ALP׫C{HK�_SCT��F_e�F_o�����FS�J�j�CHA��1��9I�s�8RS�D_!聂��恩�_�Tg�7�� �i�EM,��0Mf�T&� @��&�#�DIAG~��RAILACN���M�0�"��1����L��{�PRB�S&   ��C4�&��	��FUNC�"N��RIN�0 "$��7h�� S_��(@���`�0��`A��C#BL� u�A�����DAp�a���LDܐð�����2j��TI%���@�$CE_R�IAA��AF�Pb=�>#��D%T2� 1C��a�;�OIp��DF_Lc�X��@��LML�FA��HRgDYO���RG��HZ 7����%MULSE� �����k$JۺJ�����FAN_ALML�V�1WRN5H�ARDr��Fk2$SHADOW|� �a��O2s�0N�r�J�Y_}���AU- R+~�TO_SBR����3���:e�6�?�3M/PINF@{��4���3REG�N1D�G�6CV��s
�F�LW��m�DAL_N�:�����C	д���a�U�$�3$Y_Bґ u�_��z��� �/�EaG��ð�AAR�������2�G�<�A�XE��ROB��R�ED��WR��c�_�M��SY`��Ae�VSWWRI���FE��STՀ����d��E"g�)��D-�{2���BUP��\V��D��O�TO�1)���AR�Y���R���bנF�IE���$LIN]K�!GTH�R�T_RS���E��Q�XYZ��Z5�VOFF���R�R�X�OB��,8d����9cFI��Rg���4��,��_J$�F�@貿S��q0kTu[6�� 1�w �a�"�bCԀ+��DU�¤F7�TU�R0X#�e�Q�2X$P�ЩgFL�Pd��㐗@p�UXZ8���� W1�)�KʠM�䂤F9���ӓO�RQ���fZW30�B�OPd�,��t��8��A�tOVE�q_BM���q^C�udC�ujB��v�wL�wg��tAN=�Q�qD!`A�q�� =�}��q�u�q���dC���"���ERϡj	B�E��T�ńAs�@�UeX��W����AX��F����N� �R��+��!+�� *� `*��`*��`*�Rp*�xp*�1�p*�� '��  7�� G�� W�� g��  w�� ��� ��� ��đ޸�DEBU=�$�8D3�h����RAB�������sV��<� 
��i�`A��-� �������a���a�� �a��Rq��xqJ$�`D"\�R9cLABOb�u9�F�GRO��b=<��B_���AT� I`�0`����u���1��ANDfp�ຄ���U���1ٷ ���0�Q�0������PNT$0M?�SERVE�y@�� $%`dAu�!9�PO��[0ЍP�@�o@*�c�x@� � $]�TRQ"�2
\��Bf��j�D"�2�{�" � _ �� l"T�c6ER)Rub�I��VO`Z�N��TOQY�V�L�@P)�1R�Ƅ G;�%�Q��2 [�T0e�� ,h7�ř��]�RA#�? 2� d@��ӹ�r� �Y@�$�p�t ��OC|�f��  �˟COUNTUQ�F�ZN_CFGe��# 4B�F��Tf4;�~�\� �
�ӭ�uC� ���M: �"`A`��U��q: �FA1 d�?&�X�@=����H_B�A<����AP���o@HEL@���� 5�`B_B;AS�3RSRF E�CSg�!��1
ת��2��3��4��5*��6��7��8
ל�ROO�йP�PNLdA�cABH�� ��ACK��INn�T��GB$Uq0� +\��_PU��@0��OUJ�PHH���, u���TPFWD_KcAR��@��REG�� P�P�]QUEJRO�p�`2r>0o1I0�����P����6�QSEM��O��� �A�STYk�SO: �4DIw�E����r!_TM7CMA�NRQ��PEND��t$KEYSWITCH���� �HE�`BEATM6W3PE�@LE��]�|� U��F>��S~�DO_HOMB �O>�_�EF��PR�>a9B�ABPx�COx�!��#�OV_M�b<[0# IOCM�d'feQъ�HKxAG� D�QG��Ue2�M�����cFO;RCCWAR�"�����OM�@ � Q@r�:#�0UHSP�@U1&2&&3&&4�AT��s�O��L"�,ҞHUNLO��c4�j$EDt1  �SNPX_AS�҇� 0+@ @��W1�$SIZ�1$V�A���MULTI�PL��#! A!?� � $��� HNS`�BS�ӂAC����&FRIF�n�S���)R� NF�ODBU$P���%B3=9�G�Ѫ�y@� x6��SI��TE3s�r.�cSGL�1T�R$p�&�П3a�P�0ST�MT1q�3P�@5VByW�p�4SHOW�5n��SV��_G��;� Rp$PCi�oЬ���FB�PHS�P' Av�Eo@VD|�0vC�� ���A00޴RB% ZG/ �ZG9 ZGC ZG5XI6�XI7XI8XI9XIAXIBXI ZG3�[F8PBZGFXH��XdI1qIU1~I1�I1�I1�IU1�I1�I1�I1�IU1�I1�I1 Y1YU1Y2WI2dI2qI2~I2�I2�I�`�XP�IQp�X�I2�I2�IU2�I2 Y2Y2Y��p�hdI3qI3~I3��I3�I3�I3�I3��I3�I3�I3�I3��I3 Y3Y3Y4�WI4dI4qI4~I4��I4�I4�I4�I4��I4�I4�I4�I4��I4 Y4Y4Y5��y5dI5qI5~I5��I5�I5�I5�I5��I5�I5�I5�I5��I5 Y5Y5Y6��y6dI6qI6~I6��I6�I6�I6�I6��I6�I6�I6�I6��I6 Y6Y6Y7��y7dI7qI7~I7��I7�I7�I7�I7��I7�I7�I7�I7*�I7 Y7Y7T��VP� Uc�� l�נ��
>A820�����RCM2���MT�R��|���Q_��R-��ń�����[�YSL�1�� � �%^2��-4��'4��-Y�BVA�LU�Ձ���)���F�J�ID_L���H�I��I��LE_������$OE�S�Ab�� h �7�VE_BLCK�¡1'�D_CPU7ɩ 7ɝ ������E���R � � PW��>�E 6��LA�1Saѝ������RUN_FLG�Ŝ������ ����������H���ЧĽ}�TBC2���/ � _ B��� �br� W?�eTD	C����X��3fՆS�THe�����R�>�k�ESERVEX��e��3�2 �d���� �X -$��LENX��e��Ѕ�RA��3�LO�W_7�d�1��Ҵ2& �MO/�s%S80t�I��"�ޱH����]��DEm�41LACE��2�CCr#"�_�MA� l��|��T#CV����|�T��� ����0Bk�)A�|�)AIJ��%EM7���J���B@k�X�|���2�p �0:@q�j�x JK��VKX������f��J0����JJ��;JJ��AAL����(������4��5�Ӵ �N1�� ����L�F�_�1� 	�CF�"� `�GRO�U���1�AN6�C��#\ REQUIR��4EBU�#��8�7$Tm�2���p|ё %�� \�/APPR� CA��
$OPEN�C'LOS<�Sv��	rk�
��&� �<��MhЫ���v"/_M	G�9CD@�C ܺ�DBRKBNO�LDB�0RTMO!_7ӈr3J��P��������������6��1�@� 9$��� � ���'��-#PATH)'B!8#B!��>#� � �@�1S�CA���8INF��UCL�]1� C2@UM�(Y"��#�"������*���*��� PA�YLOA�J2L�ڠR_AN`�3L���9
1�)1CR_�F2LSHi2D4L�O4�!H7�#V7�#ACRL_�%�0�'��$��H���$H�C�2FLEX�:�J#�� P�4��F߭߿���0��� :����|�HG_D�����|���'�F1 _A�E�G6�H�Z�l�~����BE�������� ����*��X�T,�C� ���@�XK�]�o�^Av�	T&g�QX>�?��4T X���eoX�������� ����������	-	:"J@� �/�M0_q~�۠AT�F��6�ELHP���s�Jڗ � JEoCTR�!�ATN���v|HAND_VB�q�1��$� $:`�F2Cx���SW�5�� $$M,00�_Y�ni��P\����A��� 3�����<AM��_A�mA|��NP�_D*mD|P\ G��E�CSTaM�nM�NDY��� C����0 ��>7_A>7Y1�'��d�@i`�P��������"Qs$�� O�4D'"r�J���OASYMl%A�� Bl&��@�-Y1�/_� }8� �$��� ��/�/�/�/3J	<�:;��1�:9�D_VI��x���V_UNI�ӝ��cF1J����� ��Y<��p5Ǵ�y=6�@�9��?�?>�wc�4��3=��$� ASS  ���s��  ��{�h�VER�SIONp��~��
��IRT�U<�qσ�AAVM_WRK 2 ��� ?0  �5z���r����� �A	8�)�L�{����:�w�^�|�(ܛݧ�7�����������BSP�OS� 1���? <��A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� ������� #5GYk}�� �����//1/�C/U/ⰑAXLM�T��X#�%�  �dj$INs/�!i$P�RE_EXE�( � �&)0�q��������LARMRECO�V �ɥ"
�L�MDG �����[/LM_IF �ˆ!X/c?u?�? �?�:Q?�?�?�? OM, 
0�8O�4��cOuO�O�O�NGT�OL  ���A�   �O�K��PP�)�O ; �?6_,_>_P_{�  $BR_�_w�o_�_�_�_ �_�_o�_'oo7o]o�!��O�o�o�o�o�o �o�o+=Oa��PPLICATf��?��� �%@�Handl�ingTool ��u 
V8.3�0P/33�@lt���
8834�0�slu

�F0�q�z{�
2�026�tlu���_�7D�C3�pJ  �sN�onelx� �FRA���p���B�TIV�%��s�#��UTOM�OD� E�)P_CHGAPON�������ҀOUPLE�D 1��� ���"�4�uz_CU�REQ 1�� ) � >�>�*ސ�p4��!��x�~�� ��u��H�m����HTTHKY����w���7��� �%�C�I�[�m���� ����ǯٯ3����!� ?�E�W�i�{������� ÿտ/�����;�A� S�e�wωϛϭϿ��� +�����7�=�O�a� s߅ߗߩ߻���'��� ��3�9�K�]�o�� ������#������ /�5�G�Y�k�}����� ��������+1 CUgy���� ��	'-?Q cu����/� �/#/)/;/M/_/q/ �/�/�/�/?�/�/? ?%?7?I?[?m??���P�TO�@����DO?_CLEAN܏���CNM  �K >�aOsO�O�O�O�D�DSPDRYRLO̅HI��=M@NO _'_9_K_]_o_�_�_��_�_�_�_�_J�MA�X�p�4�1���aX��4"��"���PLU�GG���7���PRUC�@B;@?K_��_ebOjb�O��SEGFӀK�o�g�a;O MO'9K]�o�aLAP�O~Ǔ�� �����/�A�S��e�w���΃TOTA�L-fVi΃USENU�`�� ��䏺��P�RGDISPM+MC�`{qC�aa�@@}r��O�@f��e��_STRIN�G 1	ˋ
��MĀS��
~`�_ITEM1j�  n���������� Ο�����(�:�L� ^�p���������ʯܯ�I/O SI�GNALd�T�ryout Mo{dek�Inp��Simulate�do�Out.��OVERR�@ �= 100n�I?n cycl"�o��Prog Ab�or8�o��St�atusm�	Heartbeati��MH Faul<����Aler��� ݿ���%�7�I�[�m�� �3f��1 x�����������*� <�N�`�r߄ߖߨߺ�����������WOR�`f�L���&�t�� ������������ (�:�L�^�p�����������POd����� d���%7I[m ��������!3EWi��DEV������ ��//'/9/K/]/ o/�/�/�/�/�/�/�/|�/?PALT�� 81d�?`?r?�?�?�? �?�?�?�?OO&O8O�JO\OnO�O�O�O&?GRI`f��AP?�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o6oHo�OR�̀a�O Zo�o�o�o�o�o &8J\n�������noPREG<>%��o�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~���~��$ARG_L��D ?	����ӑ� � 	$�	[�]����Ɛ�SBN_CONF�IG 
ӛ&��%� �CII_S�AVE  ��E�<�ƐTCELL�SETUP �Ӛ%  OME_�IO��%MO�V_H������RE�P�l���UTOB�ACKt�0��FRA:\� ����_�'`����=�� J� 	������ͿĿ8ֿ�6����	�1� C�U�g�yϋ��Ϸ� ��������ߜ�5�G� Y�k�}ߏߡ�,����� �������C�U�g��y����a�  �)�_�_\ATB�CKCTL.TM�P DATE.D�;<��	��-�?��IKNI;0p�8��?MESSAGT�^��_�ېi�ODE_D ��W�8�H���O�����PAUS��!�~ӛ ((O֒ ��
��*N<r `��������"����TSK � ��=�C�	�UP3DT��\�d����XWZD_ENB8\�4��STA[�ӑ܍őXIS&�UN�T 2ӕ`� �� 	 ����0@�n���b{N��Q7���`�`'$7�  /L/^. "�YK����ď` �Ď}��=/�/a/�/��/�MET�`2��P�/?�/<?�)S�CRDCFG 1�C`��\�\�1?�?�?�?�?�?�?6��QX��??O QOcOuO�O�O O�O$O �O�O__)_;_�O�O���GR����zS���NA��қ	��wV_EDZ�1�e9� 
 �%=-��EDT-h_ʪ��_o�`/A���-(��_�	�������_�o  ���e2 �oɫko�o�6k�o! hozo�o�c3Y�o ��o�n��4F�j�c4%��r���n�N��� ����6��c5 �a�>����n���̏ޏt���c6��-�
� Q��n�Q�����@�Ο�c7����֯��n��@�d�v�����c8U��_����0
 }~�� 0�B�ؿf��c9!ϑ�nϵ� }Jϵ������2φaCR�oį9� K���������n����zP�PNO_DEL��_xRGE_UNU�SE�_vTIGAL�LOW 1�Y�~�(*SYS�TEM* 3	$SERV_GR�R� 69���REGB�q$d� <9�NUMg�<��z�PMU�� 5�LAY�  <PMPAL[�>��CYC10�����������ULSU`��{�����D�L�~N�BOXORIk��CUR_;�z�PoMCNV��;��10���T4DL!I�%9�[���ߨ ��'9K]o�R�zPLAL_OU�T Dcc�QW?D_ABOR��	���ITR_RTN���Y� NONS�8� �CE__RIA_I��5<F_1��B� =[_PARA�MGP 1�w`_���^�Cp  .� U� � � � U� � � � �� � � �  D5`D$3!g-կ<$�H$�T$�W DX � X Y"� B�D1� 9X �@� 6?� <HE��ONFIy���!�G_P��1� �e�U??0?B?�T?f?x?�?�!KPA�USX�1�UR ,Z��?�?�?�?�? OOOTO>OxObO�O��O�O�O�O�O_�2O�_ey�PCO�LLECT__0�Y5auGWEN��I��cR QNDEOS��W��12�34567890��W�S�u�_�Vy
 H�y)�_#oS� �_ohoT�AoSo�owo �o�o�o�o�o�o< +�Oas�� ������\�'��9�K���o��VQ�2�W[ � t�VIOG �YcQyH`&�8�J�\��TR�K2؍(��
��j��  ����%퉯_MOR҂!� x+ �'� 	 � 5�#�Y�G�}�k����"Ӂ"��2?�!�!H3 ҡ�Kڤ��$�R_#*_	���C�4  AS yC  �x�A3!z  �BC!�PB/!�PC�  @*���^�:d�
�IPS�$���T��FP?ROG %�*6���8��I����&R�ҴKEY_TBL�  )VR� ��	
�� �!"#$%&'()*+,-./�W�:;<=>?@A�BC��GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~�������������������������������������������������������������������������������͓���������������������������������耇����������������������1��LCKۼ3����STA�д_A+UT��O(��U��INDtTD�FQR_3T1_�Q�T2��7�$����XC� 2�����P8
SO�NY XC-56�������@����u� ��А;�HR5��cT�0�B�7T�f�Af!frꬿ���� ���� ���5�G�"�k�}�X� �������������ǼTRL��LET�EG��T_SCREEN �*�kcsc:U�$MMENU 1�&�)  < ���y��Ã �=&sJ\ �������'/ �/]/4/F/l/�/|/ �/�/�/�/?�/�/ ? Y?0?B?�?f?x?�?�? �?�?O�?�?COO,O yOPObO�O�O�O�O�O �O�O-___<_u_L_ ^_�_�_�_�_�_�_�_ )o oo_o6oHo�olo ~o�o�o�o�o�o�o I 2X�hz����� _MANUAL�ߕ�DB��L�+�DBG_ERR�L��'�� ��\�n����N_UMLIMK��d �p�DBPXW�ORK 1(��I�ޏ����&�ŽD�BTB_@ )��������qD�B_AWAY��_�GCP  �=�9װ�~�_AL��D߄z��Y��M � �_n)� 1*����
͏����6�6@�_M{�ISAЉ��@B�P�ONTIM6J� ��p�ƙ�
�ۓMOTNE�ND߿ڔRECO�RD 10}� y�>�?�G�O�� ��?���2�D�V�h��� p������*�߿�� ����9Ϩ�]�̿�ϓ� �Ϸ�R���J���n�#� 5�G�Y���}��ϡ�� ��������j���C� ��g�y������0� ��T�	��-�?���c� ��\����������P� ����;��_q� ����(�L %�4[��� ��^t�l!/� E/W/i/{//�//�/�2/�/�/??�/z�TOLERENC��sB�В��L����CSS_CNST�CY 116� 	 ?Β�?�?�?�? �?�?�?OO&O8OJO `OnO�O�O�O�O�O�O�c4DEVICE ;126� b�*_ ?_Q_c_u_�_�_�_�_��_�_?�d3HNDG�D 36�Cz��^LS 24] �__oqo�o�o�o�o�o��_e2PARAM C5�B��t�dc4�SLAVE 6�6�e_CFG �7��gdMC�:\e0L%04dO.CSV�o��c|l�r�"A �sCH�p�&a&��n��w��f�r����À�JP�>��\_C�RC_OUT �8U����oEpSG�N 9U�Ƣ���\�16-O�CT-22 14�:21�p�0�2��4��9V UBu1�݁�nހ���o��Im���P�uG��@uV�ERSION ���V3.5�.11E�EFLO�GIC 1:ݫ 	6��|�C����^�PROG_E�NB����͢��UL�S{� ��^�_A�CCLIM|���Xs��WRSTJN[���ţ�^��MO��¡Zr,�INIT ;ݪs5᡻ *�OPT$p �?	i�B�
 	�R575�c��7�4��6��7��50��R�Ƣ2��6��X�>y�TO  ���t?�Y�VP�DEX��d���@W�PAT�H A��A\�E�����7;IAG_�GRP 2@�k�,�"	 E��  F?h F�x E?`�D���û��V1"�ü��XT0K�9�Cf�py�p�Y�dC�pqߪB�i�ù�mp4m5 78�90123456���;����  �A�ffA�=q�AةpхAʯ�HAĩp����~���A��Mk,���@��tp�p���W0A�T0T0�pBA4ü Qô���
����(�A�A��
=A�L����A��
A�Q��A��������e�����e� Pe��:��{A�d������dѩp�������A�������́�r߄ߖߨߺ�@�E�G�A@�p:�R�A5d�/��)��#
P�d�l�������"�4�F�@�Pz�A�J��c�?��9p��A3\)A,��A&����0���Ю�����@�cP�]�W�AW�P�J��UC��<d�4�-d�%G��(�:�L�^� @���$HZ�� .|����bt � 2Vh�x m�����[���s������=�
==�G=��>�Ĝ���7���8��b��7�7�%�@wʏ\"&�p�.%���@�Ah�p9 A���<i��<x�n;=R�=s���=x<�=�{~Z�;��%�<'�'�~ �?�+ƨC�  <w(�U� 4"w����&����%ùf��@?Œ?� ?@?R?g��$^?�?"?��?�?�?�?�?�?)�7L?S�FB$��/"Eͽ�>OG�ΐԬq��sD�5L4�x�CA��Gb�@tφ���-_7_�C���_;�/_�NED � E�  Eh� D[PbRD_¿�_��8�?�p(�ج�Q�
'���Y�Q4����3�P����Q���ѪC=��D"	�q<�{_�_w_Do�K:o@bù�Y�7m�)6;�T�*�/9B�P o�o
o�o�o�o�o�o�ĿDICT_CO�NFIG ���Yt؃e�g��ԱSTBF_TTS�
ęVs3����
�iv[�MAU����Y�MSW_C5F*pB�  �Q��OCVIEW}pC�}���6�
�� .�@�R�d�w����� ��ȏڏ�{��"�4� F�X�j���������ğ ֟������0�B�T� f�x��������ү� �����,�>�P�b�t� �������ο��� ��(�:�L�^�pς��|KRC�sDJ�r!� �κ�������7�&��[�otSBL_FA?ULT E���x>u�GPMSK_w���pTDIAG �F.y�q�IU�D1: 6789?012345��;x�MP�o!�3�E�W�i� {������������`��/�A��( W!��J�"
��vTR'ECP����
���� �M�(:L^ p�������  $6]�o�l���UMP_OPTIcON_p�ގTR�rt`s���PME^u��Y_TEMP � È�3B��pp �A  �UN�I�pau!�vYN_?BRK G�y���EMGDI_STaA%�1!G%NCS#1H�{ �K��9�/_}dd�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO��O�O�O�O �I�!�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo �JO�o�o�o�o�O�o �o+=Oas �������� �'�9�K�]�wo���� �����oۏ����#� 5�G�Y�k�}������� şן�����1�C� U�o�]�������ɏ�� ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�g�y��� �ϧ�]�ӯ������ %�7�I�[�m�ߑߣ� �����������!�3� E�_�q�{������ ��������/�A�S� e�w������������� ��+=Oi�s �������� '9K]o�� ������/#/ 5/G/ak/}/�/�/� �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OY/KO uO�O�O�/�/�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oQOcOmoo�o�o �O�o�o�o�o!3 EWi{���� �����/��o[o e�w������o��я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�S�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�K� 9�g�yϋϥ������� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�C�U�_�q�� 9�Ϲ��������� %�7�I�[�m������ ����������!;� M�Wi{���� ���/AS ew������ �//+/EO/a/s/ �/��/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O =/GOYOkO}O�/�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo5O'oQoco uo�O�O�o�o�o�o�o );M_q� �������� -o?oI�[�m���o�� ��Ǐُ����!�3� E�W�i�{�������ß ՟������7�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �/�9�K�]�oω��� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ���������'��C� U�g��w������� ����	��-�?�Q�c� u��������������� �1�;M_�� ������ %7I[m�� �����)3/ E/W/i/��/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?O!/+O=OOOaO{/ �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_O#o 5oGoYosOeo�o�o�o �o�o�o�o1C Ugy����� ��o�-�?�Q�ko }o��������Ϗ�� ��)�;�M�_�q��� ������˟ݟ�	�� %�7�I�[�u������ ��ǯٯ����!�3� E�W�i�{�������ÿ տ�a���/�A�S� m�wωϛϭϿ����� ����+�=�O�a�s� �ߗߩ߻�������� �'�9�K�e�o��� ������������#� 5�G�Y�k�}������� ���������1C ]�Sy����� ��	-?Qc u��������� �$ENETM�ODE 1I^��  
  (/:+
 �RROR_PRO/G %*%}/��)X%TABLE  +h�/�/�/��'X"SEV_NU�M &"  ��!!0X!_AU�TO_ENB  qD%#U$_NO21� J+9!2�  *�u0�u0�u0�u0(0+t0�?�?�?N4HIS3
 �G;_ALM 1K.+ �u< +�?/OAOSOeOwO�O�?_2T0  �+s1:"�J
 TC�P_VER !�*!u/�O$EXTLOG_REQ�6s�E9 SSIZ)_�TSTKFYc5��RTOL  �
Dz�2�A T_BWD�@�P<6ܯQ8W_DI�Q L^G48$
?"�VSTEP�_�_
 >�POP_DOh_!�FDR_GRP s1M)B1d 	�O�fo: W`�������glp�w�qŗ��I ����f�Wc�o�mW`C}�X�B��FCd���A��B�ځ�B�;��mB)���A��BH��
A���A���m�o3WB�{f��p/V!�A.�>�Β�� 
 E��q �b�pr�wN��B��8�#�\��m`�}dC��N��B��{���m@UUT��UTF�Ϗj��s����m�OHcEP�]��O��#M���*�KA����m?�F��:�6:N�r�9-��z��m��+�����m��u(�<!����z��;�+FEATUROE N^�P>!�Handl�ingTool �� mpBo�English �Dictiona�ry�
PR�4D Stڐa�rd�  ox,� Analo�g I/O�  �ct\b+�gle� Shift� � !*�uto S�oftware �Update  �fd -c�mat�ic Backu�p�IF O���ground �Editސ�g �R6Came�ra3�F7�Par�t��nrRndIym���pshi���ommon ca�lib U���n�����Monito�r�CalM�t�r�Reliab�L��RINT�Data Acq�uis�Z�ϠC�iagnos��0�<��almC�ocum�ent View�e�\���C�ual� Check S�afety��  �- B�Enhan�ced Us��Fyr���8 R5��xt. DIO 6�fin� (�@ϲwend��Err�=Lm� D p^��Z��s	�EN�r.��հ �P�rds�FCTN MeKnu��v8���m��FTP In'�f�acN�=�G��p �Mask Exc���gǱisp��H�T^�Proxy �Sv��  VLO�Aאigh-Sp�e��Skiݤ e�f.>�Hf�ٰmm�unic��ons��
!
��ur�E�'�7�rt F�4�a�conne�ct 2;�Inc=r`�stru����� SpKAR�EL Cmd. �L��ua��OAD�*�=�Run-TiNưEnv� �D;�^(�el +��s���S/W�.{�License���
����ogBo�ok(Syste�m)蔭�JM�ACROs,��/�OffseS�Z�M�Hٰp��� j73�ΰMMR��l�3�5.f��echS�top��t�R� 7ize*�Mi��O� 2�7�x��0���n�miz��odM�witch����a�.�� v���O7ptm��49����fil��ORD���0�g�� 849~6�ulti-T�������CPC�M fun,��.sv�oO����� �^�5�Regiҷ�r��	�!2�ri���F�  H59�k�1�Num Se�l*�  74 H|��İ Adju����adin��O� y,[���tatub��\У�������R�DM Robot���scove� ��d em(�ٱn�� SW��Servoٰs�ꒄ�?SNPX b���1��g P�Libr<���1�ڐq 9� ɰ.30g �o��tE�ssag�� f��@ �e����"g��/I�_�
�I�TMIL�IB���� P Firmn���^�FAcc����0���T�PTX���510.� eln�����x����H573��rquM�imul�a��� 2�ToMuz�Paxѩ1� �T��6���&��ev�.��IUSBg po����iP�}a�� 0\sy nexcept��|3 <� \h51 �����oduV #��9��Q�VN�k"6PCVL{&�^�}$SP CSUI��d���+XC��a�uҠWeb Pl���t? �#S��\" 	2�������S�&ުz�V?8Gridplay��&� ���8�-iRb".� �@ � R-2000�iC/165¦ �d+�+�larm �Cause/1 e�d�<0:�Asciyi����Load��V4�3Upl�0�_�CycL�c�m�or�i����FRA[�a�m�) tdt��NgRTLi�3Onݐ�e Helݨ 5�42*�PC`ρ�4��`�]�1trߵ4�8��ROS Et�hv�t[���10�\ҠiR}$2D ;PkߵDER>1�E����of�A��ΰ�FIm��F�� z���64MB DRA�Mު�@:�9RFRO<A[�Cell3� �����shrQ
��ZcЛ��ÍUk�p� p�ide�WtyL�sL��|0\z�!Ctd���.��@"EmaiF��li���+�\��� R0�qZ$Gig�E�N�4OL�@Sup"��b�W3oa�~�cro������4���QM��Fauesat�A>�j�� miH9.dVirt��W��0{&ImM�+T����}$Ko�l Buir��n�յ'APL�&4��MyV6� "�0�*�CGP�l���{RuG�'p�{SBUW��RQ�)K�&cm\ :��z��fX�)O�v�v�(TA�&spoҠ�-�B�&��
 I�\E �P�+�CB'fg-x��&"  �E��sv�b��vv�3���S_k��TO;-�E�H�f6.
�E�vf�x_z�)�V��tr >�)�hZ%.�F�&  � ��r���*�G�&�� �њr����H��Р^JzCTIAc�pw�4�LN�1�Mr�"C #[��g�"�M�$-�P2�~T�@�����vxui�-�SD�&�S�&�*4�W���2.pc�)VGF���fxwʪVP2AU \fx���N��if�u���"inVPB���)���s�D��*�a<�s�F�5 M��zs�I��c�{&�Traİ��U,p  ��<��2��<RDp	�N��HY�<��p��-��H����Øp)����y �ϭ����ħϞ��rд����í�4+���'9Ly���ӎ��yߞ9ӫ�c3�U���B�O�q�u�y�kߍӍSy*�ߞ��\Yy����k��W���ӄ�Yyx����:�	�ߞ�����5�o��e/�Q��,y�K�m��g�^~���us�2��A��������F�������y�)���|��<��1�m�.�+�M�Ϗ�8G�i�7n��c���1�� <����W������7�{����6��Z������uk<��[�|�!�3�?�ϔ��iB\�g���_��{�x@.��wrs�t���B�� H#68��@H)xT@J�EENDI?N��tql[}
_��w�P�TQ y(��I) "���PA���T�/��'85/A#bs;/ �C/U/�,q�/B�Gp`�/�#��/�"36��5�R ?!2epai?5!:/Y4W���%INTo?e?_.q�?�4)��?�2pa2g��?�F O�?A�a�d6?��t ZUD2�gunOOqC533�R?�D�0u�O�/�Mcam���OO�LNT� ?��P_�Ĕ�0_QR7�L_�Cfi._H?_,_�f'R50�_�SAF�-F�_�7�w.v�o��_�_8�/�dM� Cbo���o�bv9rEo��paa�oaDx�@�osF-AS"-sS�p'Is(�PC�esXPL�O�tlo�_�ut\a�Oh%a9fvh%- B��/�����C�$��sr�p�?@_�?`w�}�bA�����h�`��]T�<ˏ�sgch�o2s�t��CG\s;��u1s�?���Sg�/�gG J����GDǟri$"�o�gdiʏ�!�fd���?h%J364S��Tut�o�O �?s����F�_��� �E�0���D`!�)�`NO4E�O�i$II���iwjOl�ž��>�?*�lb
��V��vjr/��
���7���2��_�?zG7\2O�E G��Ϲ?���1� ޯ&��_d�oi�8��c��50�>�x�Ͻ�"L�o�h%����dj9��﴿ƿؿ�c� u9p9�C� j9{�E�2�L��Ek,B串 ����oS_e_�&/���O}�j94JϬ�duZ��U��=d;������8���r7�Dh�u���;]m AT��������f�a���M����P��-4r V��O"3 #S�dwc�P��in�`�a�?& �HTuRef���I
�?hc�g�r"���q.JG"�er�M/��/ �/LRA�^��uH71�/�tC9K�/<eTXP/?i�9k1/m5k.f��3riR�eHG�/ƪ/ cr�NHG�Rf?L�iY�7�hOuX��H\mO��oρ� ;H��DD@�O��*�<��:I�?�?��d�R�_ 3hd�ghgOO��_���gmh�_h�m ��XO�o|O�O�o�O\/$�o0�f�gm�o`���`e۠;iov���yt��"��uR60���#tmo_�3#1��fdr,�op7��_����lp�>oh��冬~� ߏ�dgts���&dޏ�/�o�o
��J?<�vrF���v.�R���Ɵpld�5�6�%4�0/���re�eK�m�XP)�KCO*O|%56?�OZ�` o~����E$io��0��jߠ���l ����3OR��LOFvod��_IF��$�� ߪ�dDߦX!B� Uce��ft�4 ���(M�O�5)e?Ƕ/���1?Q�D�uk�'�|� ���`�boto�����-���6�p�eS ��on*���^�lB'�����Տ_�q�_�rdk��4f��C(ҿȿ ¯ԯ������̟��𒜩��
I��5s71��t�adi3f9Tar��l�ofk0�������vPa�@�� PJ��|*`��������et�&4epg���ed��� E�5�RI � H552n� 747�21�p�WelR78��,� �0ETX�J614���ATUP  wwmfh 545�p��"6�pk�V�CAM  7\a�wCRI@ EwD" G UIF)�!28  j�C�NREM�`�63��a�SCH  �4C DOCV�� CSUi�!0� D sEIO�CE�54�#R�694 we!!ES�ET=S#!3!�a 7�3!fanuM�ASK��PRXY�_"7� �0�'OCO��"3=P[�<#"�ER J�" x7�!!J774#!;39�  Eq�G1��LCH 0#OP;LG%J5000#oMHCR)%PS�1.7#MCS 4D"�0�4 O#J55 [#MgDSWe!Y1MD#1�s#OP#1#MPR$07�0w"0�#�  Σ#PCMX �#R0 A�#� &�00�#� 0( �&0�$50( �#�PRS� 3J69\03FRD@ 02�RMCNy�ndM��93 SwNBAA�800�@�HLB  "Lo��SM�A0 (W�w"4 onit#!2�  II)�TC< [#TMILe �B��`0"K3�@TP�A� �QTXa�t�\j�@EL�BM25�0`0/D8��$78n�mon�195d vSD95\FUEC 0OP� UFR@ ��;!�C@ \�@;!O�0p�t"VIP�@#� I:�@0�!CSX� �#�WEB �#HTT. \stB24 �#�CG�Q#IG�Qtwopm�PPGS!�f�PRC�@SH7�$��w!6( �8��!�[�R RBB- Ci��B01rogw!#IF#"098-!!` ��@�A64�(AaN�VD�!Ld�1h 6a6�8( c�`d SR7^c!te.p� 0ka�ч@�bc`� CLI�$0?�sb$c9G MSp�"5a�` - A� wSTY�@al �@�CTO �CJNN�0J98�ORSp�0G��b�g J�`�OL�1Abn: S�ENDu�to�!L��Q���@*r#SLM�� 8�"FVR� M�CHN0CSW!SPcBVP�� PL� �ds �qV$0�cCC�G $p�aCR�0
�Np�QB� 87.f:�QK� j70*`�p��0'3CSqToo��CTQ���qTB$�P�N��@n;pq�C�@�Q#�� �p, #�p ��. %�$07#%�� `8D#TC� QSQ"TE� [#m� �tTE� gt"m�P�T�TF�Q[����@�#C�TG�Q�"���@�#C3TH `�TTI�@#�CT'Qeqs�PCTM�@SC�$0gS�^�0bodyqP�@�  ��� �1� d��q�a�us�a9��P[�qW4 `@06; GF `8��V@VP2@ 623�R i��@j?�g� `n��g�B `" g�D� `��g�FX mna�"PVPI��+ G V��!#V	`  23ƱRVK�@Np�@CV��Q31�934.��vo R�er�ne땗����i$��r���h��0�A���37� �<�"�\srv�����b�3b�- S�r�B"0���A�J�935땿B�5 (S�O���g ��1�1�R|�j9�3땷b��EN�5��� awm�SK� Lib��� ���������@	 �"|�h�h�#땼�b�wmsk�n�E����q���py&E�  ���!�0�2�t Fuïբ6xۯm��uji-�	I&���8k��8!�� ��땼P��2�2��2�Mai'�on@��_�/r�;pڦh;Ѐ;�G��_r���!��4�\ֶORC��+�5.�� "T¦TP��,hQ�652�1��4���<�xk�����ߦ�%t�P��QrֶSB�� ch_����)��t!0�B�"̿ h�h 땇�;���c������������>�Rp� �\toֶ3���cl�W��2p�"����� �����F����b@� Qt�a�϶0t��2ܐFsȒ�76�p䵝t	� Ad���5�82��ob�|*�{�\a��FMpQ ���A�migֶ�I�or�wI�.j�rfm��Fc����@1�EYE~� Iw���R���4�,K2Х70.�E��ld,�C�� 1�PTP]���.�"AD.�F�&3 k���ask��ȍ`4����۳dֶے��ER~�7 R�ƫ/�`T�?)�e�rv榀G?Y?k?}?�?�?ӹapa��	d����rƚ4�M��te����7H9!J�d/���G�p�ac�T��<6�b`�/� QO��$vc>�",@Vg����eYW�2�5/� BJ�h�F��R5:�d���0�`��@��I_�raj��e��he}�$`��e5(Xa�@��et���1Otdj��,�_�h�\	UI�/k�jAo�FO��`^���F��r��qW65q���K z�'6ڦus W'�Cb,'��'?��n��MFR��;]�lf�ǯ�fr>֛�w�p�/�,��_U[ǀ�мn�x'_i�{��� ��O���pJ���[@�o�in7L�O�9�\^ � 1R����+mi2״h� �j��҇- f�n�t >�MA H��I  Hw5529� (Cߑ�21��leR�78�c�ߒ0AcaJ614��~�0ATUP��ܓ��545�t-f�l�6yE=�VCA�M�tFLXC�RId���o�UIFnULX �28���mo�NREu'��6q3��WQ��SCH��=Cn�DOCV�gϠwCSU1�cxr��0$�;EIO�C%tx\c��54��oQ��9T�;�ES;ET�Temo?�S��/��7S�{�MAS�K��70��PRX�Y�T�`��7��`�O�ߐOCOe�\?�3�ô`>��0{�?���|�-��on G�?�39!'ߑõ H82LCHd���@IOPLG.�tCGM?�0��GО��MHCR�Go�S��/1_�CS4�cg�m��50T��?�5x$�[���MDSWMfb.�D�����OP��oX/2L_�PR���K�����{���88�3n�CM��0iAE,��0�Ő`~�5#�\h88�+�?��D���.?���4��0D�3��o�S4�����9��,iFR�Dd�/2E/��M;CN5�H93�K�oSNBA�U"R��7HLB��SM�՛�8��T���J52�Sa�ߐTC4�\�TTMILe��P��䴝A|�TPA���T�PTX��5��TE�L�ԫ�0䴈P��8`�˳���K�95��v��95��888��wUECd�rt �GUFRd�__�Cd�;2e-�VCO4��GVIP�;��I�T;AX~�CSX������WEB4����H�TT4�ka��2T�2�M/So�G#��Q�IG��< .�IP�GS=t\rxO�RC��aߐ7�/a��16D�s@>�R7#��! ��Oq�Ҥ��P��Ҷ�;�A���KÑ�$�0 �"��4����NVDx4���#�Adap���8D���68����R�7���P��D0��a��o�bܠ. CLIƔ�l\-C���CM�S�'��4�d "�ްSTY�[�CTmOT�tl��NN����ORS4�;�1 ��7ltiΰOLS�( AE���0�T���L��6�@���9@ ��L�M4�HV o�V�R���CS��shc>�PBV4䫁/��PL�
APV��u;st>�CCG4��0�nCR�4 H5���B���K�H573���?�����\cms�#�st.~TB���! �
�7�C�ԓ�?"�Oawsh?"��I04?"��3�TCd�K�\A 4�\sl"EĤpP��� 4�C[П"Ԥ�8c��"4�(��CT�F��c��"���C[TG�73m#G䖫THd�h� �Il��K�CTC�59m�'CTM�5M����Q0��re\g�P ���12��04��h���%S��13M�CTWd�9[@_�GmFd�SE]�P2d��t+��2�ա �2d�e[ll��PBd�I����1Dd��a�1F��t;ap VPId��ÓCV�!Vq��UA���CVK�ۣCV>#�coreL���H"�Hp!�HK"�H�atc�J�H�4$�I� �IL0H�I�2��H��H+2�IL�Y4p=�H���Ie\a�I�2 Z93�I{�H�@�NZ+��H 1��K48�Z<A�Ht{�Il �Z;"�O�Fs\!�Hk"�H {"@o�F[�PZo�Z���J��Tok�РH��H�\��Il�Z��Z2�=[ng-[gToo��I�p�j(�njrob9t_�Xbt.�JL� iur�o�I��i�!���F��POz�lin�g�j��y���Y"r�^zۢ�I�p��Gea�t^j�]��Z��_je �����_��lkҠHAm,��H|��Z��A�I�  �_�  ����Gvhm�J{�sqvnj���H49\�Jz�@L�Ij749{P�Zt\jNj�@_�"g.pjmcal��0�fu�J��^zh�m-��_bg���o�\rͫ �1�H! j���;����MT "�(�Cu�zk��bgft��JlpX���GCT�"���Gfc]�˝2�6\fߟ�926�l\� Ίu�>m��;�Mul?�Q��#7\^�K���7-[˝ث��_�61Nj48�.� H- �H�@R:_�L^ziPe��K�Я�F8\}�}�����Ћ� � Rk,�t�icMoj+@OoQxsp-@�"�3�CS jv+}LB-[5 HNj+� co~�L��z���f�k˝lb�jl!l����-˜�k/�.�x��LЎ�kipJ/�Gon,�J\A��8��SK"�� ��uto�o B������kwm� �o��H�tp�ʜ n}��exH-�˝��x���a^jIlL�je�식i���a��/���rej�1�o�V�or�zR����e qT�Z[��[lclN��߭�SOžGZD���to�{+B�H6343N�`�SG/o���sg�a�Utui��;`�J��`�;�;ndm�ndiN�{/ �/�/�/�/�/�/�/?`?/?A?�?��riΪ{! -Kj950/�sn �zk]895n/��O�t �Z��ws�g�K,�>��iag�� SGJ�Ю�o�gu���KO]Ltw�>_@	J64�1�sέ{F O>ګcdHݛ��`3_��r-�V�N74�y-�3��wRINnzlly���(m^���L���sg=c�zI" #?
+�oߡ\tw/��0�.�@�"���f�_�[yr�Kmm�K}dct^��t]�+�
PRZW7CHK
k,�;;`�y<p��lK���L.N*R85j �@_j�R ���tiN�g; WJhecN�L��F����wlZ|*��dat�ʛ�g�reN��o  �STD�r7LANG�Aoc�e�`��Q�y7��R870㕼{��8 (P�ogge���!��58\�PATT�s�� �t\��c "B�@V��1�Opatd���O����������{q㕔�5B�a�p[�m�\���7�\aw��@�a��p6�����ϯ�Ogmon���d� �0�B�m�;A��\ ö�K�I�MHCR��51 H����g�\o��@��R]� H#54ۿm�<@E���p;!�����omm�$;a��R�|�N㕬0�F�C��W�P�)Ai�6�� Fƫ�{��it�x�#{ ��iai�o����De6�ev9e����72 R�@tRƜPg��adl���nt��KRB�T�tOPTN�`772'�CTK�"'�g�(䔠�)� "AZ'�;q'�q'�'tzn&�{ E'�A{ma��- Mu���ncInDP�N�������87S2��|�d��(���������#���ma{sy��y "M��0o��䃲��et����\p1�����\ ��f���lZ����lp���9���`��+ V��ail��?��䇢�䄓���zd�<�k`��7�3.f��irdg.��- i��e\ ������ S0j�021"�1W ��(�`�4�n� (i��e,"�� "���+���coKre_�I��l`F��AY��AB��@�����H�����ABIC���Par;�M�ai�������<� c\ΖITX>���  {����1��wg Jclib��ShiW�4�� t�994\�VSS�F��� tt\j9�f "O�w� t��$%ini�/��pٰ t�5G�&,� t'\vsR&x�L�%w� tamclS/+rGef.�%#� tj�%m�� t[A�&4\9z�/�,z_v�%A8�%�a�%_ol6��8l% �%end�/<!c?.?@?R5o[?m>8�6�/�dshf�/+trt�?<OAE�'F  !�G��$%��Ƙ5vi�6���6 J�92�F3��%25 	(�%�@e&�P�%k�4O dnwzF��T�&`�XEpn�&g��?� nw\n�?�,n�d�V��N;XnF j���%se�V I/�
&�q&фU��5r w�%/F� �F�_�rclR&0\pw/Y��90�Eo`/"5�Of "U//A+dp�rm�%g¨%�Xrsu/kmS�T_ L`�6/OŔpM�LO�j��nO1|h�ODnon�|YCwrpR/�l���E�<�Pe\ga��Kr�gas�o�k��f�v��4xtf�?m$ra�o�la0�omk�_�TamN6+�4�`'9K0.v�Wې�%d�@�Ft��XE sV���ДJ737�%|�*�%,P��hB 9"+��KwcfF& �I����998�vt;omzFut vV�_�	o;�YC���:8\HF&�Y/� 0��f��deb^V��$�0�zFؠ"��g���<9)\�&��9�Wr}  �su"�st�G��X ؖf� U (�fag�n�F PzFϜ�Viaf�TX����vd���w��g��HzF- OƂW CH� �$723�F���E(A�ÿտ`2蚽Wc��WsvF&3 S�W�JR6��_�RVo RV���ӊ���vt�M\et(F�XoN�o�Fr��x����+�1T�F?teR�� J58�O  {34	Wgle,�%,�j�Dq\t"��zFfwIta1lUTA�VdϜ�gw韗Mad�Wp�Oa���6d M���e�FT��90 Hv�%NT��R69�ָ����ir\ʆM�IR��ӊenʆv���F|�3��ITCP���Ta0�p���(M�M7G�eT�o \t�pʆI��YBbusJ׈�m��I�@zFȀ���F�����/��W�'g, ��4`R_(!�sw�&s_YC67\JF��Tf_����D�fw��W��4ach�g��a96_��� _샏�_rV�%� 99YA�e���$FEAT�_ADD ?	������  	�$YA// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�o�o# 5GYk}��� ������1�C� U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿�������DEMO N~�   �� *� �2�_�V�h��� ������������%�� .�[�R�d��������� ��������!*W N`������ ��&SJ\ �������� //"/O/F/X/�/|/ �/�/�/�/�/�/?? ?K?B?T?�?x?�?�? �?�?�?�?OOOGO >OPO}OtO�O�O�O�O �O�O___C_:_L_ y_p_�_�_�_�_�_�_ 	o oo?o6oHouolo ~o�o�o�o�o�o�o ;2Dqhz� ������
�7� .�@�m�d�v������� ƏЏ����3�*�<� i�`�r�������̟ ����/�&�8�e�\� n���������ȯ��� ��+�"�4�a�X�j��� ������Ŀ����'� �0�]�T�fϓϊϜ� ����������#��,� Y�P�bߏ߆ߘ߲߼� ��������(�U�L� ^���������� ����$�Q�H�Z��� ~�������������  MDV�z� �����
 I@Rv��� ���///E/</ N/{/r/�/�/�/�/�/ �/???A?8?J?w? n?�?�?�?�?�?�?O �?O=O4OFOsOjO|O �O�O�O�O�O_�O_ 9_0_B_o_f_x_�_�_ �_�_�_�_�_o5o,o >okoboto�o�o�o�o �o�o�o1(:g ^p������ � �-�$�6�c�Z�l� ��������Ə���� )� �2�_�V�h����� ��������%�� .�[�R�d�~������� ������!��*�W� N�`�z���������� ޿���&�S�J�\� vπϭϤ϶������� ��"�O�F�X�r�|� �ߠ߲��������� �K�B�T�n�x��� �����������G� >�P�j�t��������� ����C:L fp������ 	 ?6Hbl ������/� /;/2/D/^/h/�/�/ �/�/�/�/?�/
?7? .?@?Z?d?�?�?�?�? �?�?�?�?O3O*O<O VO`O�O�O�O�O�O�O �O�O_/_&_8_R_\_ �_�_�_�_�_�_�_�_ �_+o"o4oNoXo�o|o �o�o�o�o�o�o�o' 0JT�x�� �����#��,� F�P�}�t��������� ������(�B�L� y�p����������ܟ ���$�>�H�u�l� ~��������د�� � �:�D�q�h�z��� ����ݿԿ��
�� 6�@�m�d�vϣϚϬ� ���������2�<� i�`�rߟߖߨ����� �����.�8�e�\� n����������� ���*�4�a�X�j��� ������������ &0]Tf��� �����", YPb����� ���//(/U/L/ ^/�/�/�/�/�/�/�/ �/ ??$?Q?H?Z?�? ~?�?�?�?�?�?�?�? O OMODOVO�OzO�O �O�O�O�O�O�O__ I_@_R__v_�_�_�_�_�_�_m  h$o6oHoZolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ߀�߲����������  ��(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: L^p����� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p����� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺߠ��������� 	�,�>�P�b�t��� �����������(� :�L�^�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_��_�_�_�_oi�$�FEAT_DEM�OIN  d��D`�`,dINWDEX9kHa�,`�ILECOMP �O���za�Gb'ep`SET�UP2 Pze��b�  N ��amc_AP2BC�K 1Qzi G �)h�o�k%�o`}`Ae�o m�o� ��V� z�!��E��i�{� 
���.�ÏՏd����� ���*�S��w���� ��<�џ`������+� ��O�a�🅯���8� ��߯n����'�9�ȯ ]�쯁���"���F�ۿ �|�Ϡ�5�ĿB�k� ����ϳ���T���x� �߮�C���g�y�� ��,���P����߆�� ��?�Q���u���� :���^������)��� M���Z������6��� ��l���%7��[ ��� �D�h���i�`P�o }2�`*.VR`� *c�����JPC��� �FR6:�.�4/�TX`X/j/��U/�,;`%/�/�*#.FM�/�	��/�<�/<?�+STM@G?q?��]?�=+?�?�+H�?�?�7�?�?8�?EO�*GIFOOyO��5eO"O4O�O�*JPG�O�O�5�O�O�OM_F�JSW_�_� S�n_+_%
Java?Script�_�O�CS�_o�6�_�_ �%Cascad�ing Styl�e Sheets�0o� 
ARGNA�ME.DT_o��0\so1o�Q�d�o`o}�`DISP*�o �o�0�o7�e)q8�o�
TPEINS.gXMLg:\{�9�aCustom� Toolbar���iPASSWO�RD.�FRS�:\�� %P�assword ?Config@�� ���������r�� ���=�̏a�s���� &���J�\�񟀟��� �K�ڟo�������4� ɯX������#���G� ֯�}����0���׿ f������1���U�� yϋ�ϯ�>���b�t� 	ߘ�-߼�&�c��χ� ߽߫�L���p��� ��;���_��� ��$� ��H����~����7� I���m������2��� V���z���!��E�� >{
�.��d ��/�S�w �<�`�/ �+/�O/a/��// �/�/J/�/n/?�/�/ 9?�/]?�/V?�?"?�? F?�?�?|?O�?5OGO �?kO�?�OO0O�OTO �OxO�O_�OC_�Og_ y__�_,_�_�_b_�_ �_o�_�_Qo�_uoo no�o:o�o^o�o�o )�oM_�o�� 6H�l���7� �[����� ���D� ُ�z����3�ԏ i��������ßR�� v�����A�Пe�w� ���*���N�`���֦��$FILE_D�GBCK 1Q������� ( �)
�SUMMARY.�DG����MD:�3�s���Dia�g Summar�yt���
CONSLOGi�L�^��������Consol�e log����	?TPACCN�R��%:�wς�TP �Accounti�nρ�FR6:�IPKDMP.ZIP�ϯ�
���σ����Excepti�on ߱�_�MEMCHECKm�Կb�����Memor?y Data��֦�LN�)n�RI�PE�\�n����%�� Pack�et LϺ��$ySA���STAT������ߋ� %~�Status��<�	FTP����r������mmen�t TBD��� �=�)ETHERNEU���B�S������Ethern�(��figura�߇���DCSVRAF���������� verify �all٣M(=��DIFF�����/diff�PB���CHGD�1�x� X�FQ&��	28�� 5�YGD3���'/� �N/�UPDATES.m �S/��FRS:\�k/�-��Upda�tes List��/��PSRBWLOD.CM�/���"��/�/�PS_RO�BOWEL1���:GIG�ߊ?/�?�ֿGigE ��n�ostic*�ܢN��>�)�1HADOW�?�?�?5O���Shadow ?Change��٤�&8+�2NOT�I��O"O�O��N?otific��\O٥O�A��_�� 2_կ?_h_���__�_ �_Q_�_u_
oo�_@o �_dovoo�o)o�oMo �o�o�o�o<N�o r��7�[� ��&��J��W��� ���3�ȏڏi����� "�4�ÏX��|���� ��A�֟e�����0� ��T�f���������� O��s�����>�ͯ b��o���'���K�� 򿁿ϥ�:�L�ۿp� ���Ϧ�5���Y���}� ��$߳�H���l�~�� ��1�����g��ߋ� � 2���V���z�	��� ?���c���
���.���R�d�����������$FILE_� P�R� ����������M�DONLY 1Q����� 
 ��)�@_VDAEXTP.ZZZ���p�G�L6%N�O Back f�ile !��U3�M��7���� G�&�J\�� ��E�i�/ �4/�X/�e/�// �/A/�/�/w/?�/0? B?�/f?�/�?�?+?�? O?�?s?�?O�?>O�? bOtOO�O'O�O�O]O��O�O_(_��VIS�BCK����*�.VD)_s_�@F�R:\BPION\�DATA\^_R��@Vision VDt�_�O�_�_ _o_Ao�_Rowoo �o*o�o�o`o�o�o �o�oO�os�@� 8�\���'�� K�]�������4�F� ۏj����̏5�ďY� �j������B�ן� x����1���ҟg����MR2_GRP �1R���C4�  B�O�	 �
������E�� �֯�r���OHcE�P]��O��#�M��
�KA����?�&�r���:6:N�R��9-�Z��A��  v���BH��C`}dC��N��OB�{��r���xпὫ�@UUT���U����/Ϫ�>���>c��>r�а=ȫ�>�i�=���>�����:��:���:/:6?)�:��~ϗ� 2ϔ��ϸ������z�_CFG S��T  �a�s߅߾0[NO ���
F0�� ��/\R�M_CHKTYP  ���O�����������OM��_MsIN��L����v��X��SSB7�]T�� ���5�L�,�U�g���TP_DEF_OW���L�����IRCO�M�Ѝ��$GENOVRD_DO�ֹ	��THR�� �d��d��_ENB��� ��RAVCr��U�UQ �Υ m�X��|������n�� � �OU��-[��O�������8�:���x
,.  C�x ��h�������B��ϡ�����n�!�SMT'�\.���+�w�$HOSTC7�{1]K[�Y���� MCL���MI�  27�.0�1�  e}��� /*��1/C/U/g/�!/#	�anonymou�s�/�/�/�/�/? L��8;{}/j? ��?�?�?�?�?/�? OO0OS?�?�/xO�O �O�O�O?UO+?=?_ QOs?1_b_t_�_�_�? �_�_�_�_o'_]OoO Lo^opo�o�o�O�O�O _o G_$6HZ l�_������o 1o� �2�D�V�h��o �o�o���ԏ��
� �.�uR�d�v����� ��?�������*� q�����������ݏ�� ̯ޯ��I�&�8�J� \�n���ǟٟ��ȿڿ ���E�W�i�F�}�j� ���Ϡϲ��ϋ����� ��0�S�Tߛ�xߊ� �߮�����+�=�?� �s�P�b�t����� ���������'�]�o߀L�^�p�����/E�NT 1^�� sP!���  ������*��N r5~Y���� ��8�\1 �U�y���� �4/�X//|/?/�/ c/�/�/�/�/�/?�/ B??N?)?w?�?_?�? �?�?�?O�?,O�?O�bO%O�OIO�OmJQUICC0�O�O�O_�D1_�O�OV_�D�2W_3_E_�_!ROUTER�_�_�_��_!PCJOG��_�_!192�.168.0.1�0�O�CCAMPRYTGo#o!7e1@`noUfRT�_ro�o�o���NAME !~��!ROBO`o��oS_CFG 1�]�� ��Auto-st�arted��FTP��~q��� F��������9� K�]�o����&���ɏ ۏ�����Wi{X� ���o�����ğ֟�� ����0�B�e��x� ��������ү������ �Q�>���b�t����� ��q�ο����9� ��L�^�pςϔϦ�� �����%��Y�6�H� Z�l�3ϐߢߴ����� ��}��� �2�D�V�h� ��������������� 
��.�@��d�v��� ������Q����� *<������� ��������8 J\n��%�� ���EWi{} O/��/�/�/�/�/� �/??0?B?e/�/x? �?�?�?�?�?/+/=/ �?Q?>O�/bOtO�O�O �Oq?�O�O�O_'O(_ �OL_^_p_�_�_(�`_ERR _z��_�VPDUSIZW  9P^S@��T�>�UWRD ?�EuA�  guest3V�$o6oHoZolo~o�dS�CD_GROUP� 3`E| Iq�?YM �nCON��nTAS�nL��nAXP�n_E�o9P�n��RTTP_AU�TH 1a�[ �<!iPendCan�g�~@}9PJ��!KAREL:q*���}KC�����pVISI?ON SET�`E��I�!\�J�t��s�� ��������Ώ��-����dtCTRL �b�]~�9Q
`��FFF9E3�9�DFRS:D�EFAULT���FANUC W�eb Server����bvodL���'�9�K�]�o��TWR�_�`FIG c.�e�R���Q�IDL_CPU_kPC9QB�@�� BHǥMIN�Ҭ�a�GNR_I�O�Q�R9P�XɠNP�T_SIM_DO��!�STAL_oSCRN� �y��+�TPMODNT�OLY�!���RTY�8��&�9�hpENB�Y��cƣOLNK 1d�[�`������1�C�U�ͲMA�STE���&�O�SLAVE e��_˴jqO_CFG�sϦ�UOD��Ϩ�C�YCLE�Ϧļ�_?ASG 1f���Q
 W�9�K�]�o� �ߓߥ߷���������p�#�_��NUM�S��b�U
��IPCH���j�O_RTRY_CN��Z��U�O_UPD�S���U1 ������g�θ`���`ɠP_MEMBERS 2h��` $�e�>���HyɠSDT_ISOLC  ����r�\J23_D�S��q���OBP�ROC��%�JOGv�d1i��89Pd8�?�.�D��.�?�?�?OQN s��V����3W~���������>��POSRE��$��KANJI_m�K��i�pMON j�k~�9Ry���@�//�^�r��k���9%Th��p_L��I�l�kEYLO�GGIN���`�����U�$LANGUAGE ������ �!�QLeG��lq�9R��9P�x�p�  ��Z砬9P'03X�k����MC:\RSCH\00\���� N_DISP m��DAMK�SgLOCw�آDz ���A�#OGBOO�K n���9P0~��1�1�0X�9O %O7OIO[OmN�Mɱ���I��	�5Ib�5��O�O�5�2_BU�FF 1oؽ�O2A5!_�2��=_?7 Y_k_�_�_�_�_�_�_ o�_o:o1oCoUogo��o�o�o�oe4��DC�S q�= =��͏L�O-�1CU�g���bIO 1r�� ��s20� �������� 1�A�S�e�y������� ��я���	��+�=��Q�|uE�TMl�d ����Ο����� (�:�L�^�p������� ��ʯܯ� ���7��SEV��u={�TYPl���z�����!�PRS���/S��FL 1s�}����$�6�H�Z�lό~ϯ�TP� l�i�>�=NGNAM��A5��"e4UPSm0GI��\!����_LO{AD��G %u:?%PLACi�2��3�MAXUALR�MI�c�W�T���_P�R����3�R�Cp0t�9�M���3Eݼ����P 2u��� �1V	i�00���߭�1�� .�g�xU����� ���������8�J�-� n�Y���u��������� ��"F1jM _������� 	B%7xc� ������/� /P/;/t/_/�/�/�/ �/�/�/�/�/(??L? 7?p?�?e?�?�?�?�? �? O�?$OOHOZO=O�~OiO�OK�D_LDXDISA����zsMEMO_AP���E ?��
 b��I�O_"_4_F_�X_j_|_R�ISC ;1v�� ��O�_  ���_�_�Ooo@o��_C_MSTR �w:�_eSCD 1x�M�4o�o0o�o �o�o�oP; t_������ ���:�%�^�I��� m������܏Ǐ �� $��4�Z�E�~�i��� ��Ɵ���՟� �� D�/�h�S���w���¯ ���ѯ
���.��R� =�O���s�����п�� ��߿�*��N�9�r��]ϖρϺ�PoMKCFG ynm���ӿLTARM_��z
�����и���6�|>�s�METPU�Ӷ�І�viND��A�DCOLXի�c�C7MNTy� l�g` {nn��-�&���|��l�POSCF��=��PRPM�����STw�1|�[ {4@�P<#�
g� ��g�w��c���� ���������G�)� ;�}�_�q������������l�SING_C�HK  |�$M/ODAQ�}�σW���#DEV 	��Z	MC:WHOSIZE�M�P�#TASK %�Z�%$123456�789 ��!T�RIG 1~�]l�U%�\!�S
K.��S�YP�69�"EM_INF �1� �`)AT&F�V0E0X�)��E0V1&A3�&B1&D2&S0&C1S0=�)ATZ�#/
$�H'/O/�Cw/(A�/�/b/�/�/�/?  �&?���/�?3/ �?�/�?�?�/�?�?"O 4OOXO??�OA?S? e?�O�?�?_CO0_�O �?f_!_�_q_�_�_sO �_�O�O�O�O>o�Obo �_so�oK_�owo�o�o �o�_�_L�_o#o ��Yo����o $��H�/�l�~�1�� Ugy���� �2� i�V�	�z�5�������|ԟPNITOR���G ?k   	EXEC1�ê�2�3�4�5��� �7�8�9����������(� ��4���@���L���X����d���p���|���2���2��2��2��2���2Ũ2Ѩ2ݨ2��2��3��3��3�(�#R_GRP_�SV 1�� �(��@@w�Y��=�N4"⸿�������R�_Ds����P�L_NAME �!���!D�efault P�ersonali�ty (from� FD) ��RR�2�� 1�L6�(L?����	l d��nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲�����B2]���*�<�N�`�r����< ����������,�>�@P�b�t�����BJ�  �\ � �  �� � ��  A� W B��T��� �
������� g ������B��p���  CH C�H P Ez � E�� E�` E�;%��Z�*� �  E��F[�@&��T Ai� dx�H �x�	$Hxd�
dڭ�}`( d��8(xx$$y Xtd D (DDdp WwX��	X�v@XHX���/yJ�y (� !���  7%E	��Em�Xw$%XH$%P�� �/�/�/�/ �/�/??+?=?O?a?s=F�r?�?�?�?��6��E���E�A���2��� C ���?Kزd�3 �4,O:IO\OjG�0���|MTCҷ'4 ?� W%�O�O>�N  �H�O��JA  A��C��C��_�OC_9W�  � TB�LY��
��_��\�@Q�Y=�CÈ��V�`HR0� ʒP/( @7%?��a��Q?ذaر@�6��&س��2n;�	�lb	  ����p�X��U�M`��X � � ��, �rb��K�l�,K���K���2KI+�KG0_�K �U�L2o��E	O�n��6@� t�@�X@�I��b`�o�C��N����
���}v������` q�m�|�kQ�
=ô��  Hq�o~`!b���  ��a� �B����ذa�s�G��}�m��o�q��v�O��E	'� � 0��I� �  �� Q�J:�È~T�È=���l��b@|���}~�Q����RSD���yN8���  '�<��p?���b!p��b){�B��?�C�IpB  X��ذ���C�A�av �� {��	�o�Q�IB  P��8�����P��ԕرD �O���O���A�,�>�Š
�`�l�1�	 ٩�p��� p` l`:�GT  �t�?��ff{O��įV� �P����aa�!�/�K?Y)R�a4�(ذ]�Pf����a\c\dƃ�?333-d���;��x5;��0;��i;�du;?�t�<!�+}�o�ݯ��b�Sb�P?offf?��?&���T@��A=#$�@�o[,ž� x�	�&f6�ed�g�� �Hd㯸ϣ����� � ��$��H�Z�E�~߾�&eF��mߺ�i����U���y���2���E�0����y�d��� �����������?� *�܏r�8�.o�ߺ�� ��T�);ڿP b���������P��A��T �C�=�ϵ��Y}Ɂ�2������ĶC��W�C�= ��` Ca�����Ѕ�(!�`�<����bC@_;C9��BA�Q��>V{È�����Y�u�ü��
/�S���Q��hQ�A��B=�
?�h�Ä/iP���W��ÈK��B/
=�����Ɗ=�K�=��J6XK�r�#H�Y
H}���A�1�L��jLK����H:��HK��/0	bL� �2J��8H���H+UZBu�a?�/^?�? �?�?�?�?�?O�?O 9O$O]OHO�OlO�O�O �O�O�O�O�O#__G_ 2_k_V_{_�_�_�_�_ �_�_o�_1oo.ogo Ro�ovo�o�o�o�o�o 	�o-Q<u` �������� �;�&�K�q�\������Gϭ���� C��aɏ Ĉ��<��CVF������+b� ��K<c�f�� 
E�����T�ٟt�(t��_ʙh۟���������N�������3l�C�(�:�H����T�f��t�.3��}����k���q'�3�JJ�� ���گ���4�"�]%P̲Pf��������⟛�ſ���Ի� ���/��?�{?�N�u�  fUh�*ϳ� �������Ϣ�t�.��R�@��X�bߘ߆���)Z�ߺ�  ( 5�	�������B�0�f�t�  2� E%p"E[-@��N�"B�C��%@ ߏ��%������)�;��������������%n�n�%T��%��Xc
 ��!3EWi{ ��������b*[��P�I��v�$MSKCF�MAP  ��?� ^������pDONREL7  X�[���DEXCFENB�
Y�FNC���JOGOVLKIM�d��dDWKEY��%_PAN�""D�RUN�+SFSPDTYw�����SIGN��TO1MOT��D�_CE_GRP [1���[\�� �/��?&?��?Q?? u?,?j?�?b?�?�?�? O�?)O;O�?_OO�O �OLO�OpO�O�O�O_ %__I_ _m__f_�_�O�DQZ_EDI�T�$UTCOM_CFG 1�Q��_o"o
�Q_/ARC_�X���T_MN_MOD죐�$�UAP�_CPLFo�NO�CHECK ?Q W����o �o�o�o'9K ]o�����v�NO_WAIT_�L�'�W� NT�Q�Q���_ER�R�!2�Q��� A�_t�������*P��Ώ�d``OI��P��x :q�t�C+����XG��k�)�70�������8�?��4�ӏ��d�B�_PARAMJ��Q����_����s��� =��345678901��� � ��?�Q�-�]�����u�0��ϯ����������7�ODRDS�PEc�&�OFFS?ET_CAR�PKo�m�DISz�K�PE?N_FILE���!�$a�V<`OPTIO�N_IO
/!аM_PRG %Q�%$*	�ά�WO_RK ��'�� ��K�7U��h��f�(�f�	 a���f�7���M��RG_DSBL  Q�����L�RIENTTO* ��C���Z��M��UT_SIM_D�طX+M�VQ�LCT �%��R_�x$aQ�'�_PEXh`ܜ�b�RAThg d�b�r�UP )�5� � �����X������$��2�#��L6(L?}��	l d'� O�a�s������� ������'�9�K�]�@o���������H�2>� ����/ASew�N�<����� ��1CUg�yH���P��� �  �� � �U�A�  B���PB�����H��  ����U�B�p�������N�P E�z  E�� E_�` E��;(�����Z�/�~��  E��''l���@#���T�AJ(��E!Y! a!)!m!Y!u)%)!Y!(E!�%E!ڎ$�^$A! �	!E!a!�%%	-Y! Y%�-58�Z 99HU%E!�D!	$D%% E!Q481X291�%�)95 �/W#95)%91m5a!�5)/Z7��Z (�8�1a�<a1 EE	�(�Em�494X6E9=8)%E15�� |O�O �O�O�O�O�O�O__80_B_T]F�S_y_ �_�_�Vh�����_�[��͔on�_=o�Kg�]�]&�'4 � W%po�oX� g��g�o�j�A�A��c������o�o$w���tB�(~ΐ��r�|B�` q�y�$�O���1�'k�'ۆ�3�`��0���P�( @ED�D��q?�Q�C�Z7}��o  �;�	lD�	u� ����p�X�[�2���X � � ��, �W�ΐH���9H�H���H`�H^?yH�R�l����_����	�#�B#�B� C4ӄ����c��9���
=���� ������c�Bz��Βa�m�另b��s�� �q���g䟒����Ǒ�ٖ�o���e	'� � ��I� �  ��q<�=���89�K�E�@a�g� b���������E���䮟�N��  '۰��Ɓ"�B�Ղ���т6��� �  O��C�a��	ŀ~��p=�Bp��Н� ���px����D��o�޿�o��&��#��5�Ю`Q��	� ٠U�f� �U� Q�:���#�>���?�ff\o����;� �p����F��8� ��?Y
r�$�q=�(� B�PK�f����A�A���?333���Ł;�x5;���0;�i;��du;�t�<�!��y������t����r�p?fff?�x�?&���@���A#	�@�o[�	]����� �uI��wh���-��ϝ� ���������	���-� ?�*�c�u�L��������4�V�X����EjPf��^I�m ���� �$ ��W������ �9��/ /��5/ G/�z/e/�/�/�/�/��`�A��$�t�/ �C�/"?�(d��>�?��Pn?�/�?}?�m�(��W�?C�@�` CT��?�j4�j0i1A@I��!���bC@_;�C9�BA�Q�>V`.�È����Y��uü��
��?�3��Q��h�Q�A�B=?�
?h��iOJp���W�����K�B/
=����Ɗ=�=�K�=�J6X�K�r#H�Y
�H}��A�1��=L�jL�K���H:���HK��O�@	�bL �2J���8H��H+?UZBu�?F_ �OC_|_g_�_�_�_�_ �_�_�_o	oBo-ofo Qo�ouo�o�o�o�o�o �o,P;`� q������� ��L�7�p�[���� ����ȏ�ُ���6� !�Z�E�~�i�{����� ؟ß��� ��0�V�8A�z�e�Gϭ����� C�a�/�� �爓�ЯׯCVF������üKG�b0���KH�K�� 
AEp�s�9���� (�!ϳ_�h��y���<�a5�N����T�3lC���-���9�Kϰt��.3��}e�w�k����q'�3�JJ�͑��Ͽ�����(��B5P��PK�Zgt�ǿ�ߪߕ�������������$��{$�3�Z�  fU M���������`Y��7�%��=�0G�}�k���)Z����  ( 5��  ������'KY�  2 E%pnIFE[@tN�IF�B�!�!� C��0� T�@į����*H3��Tf�x��T�T�"a4��T�D=4H;
 �//*/</ N/`/r/�/�/�/�/�/��/�/GJ@2��5�I��v�$PAR�AM_MENU �?����  DE�FPULS��	�WAITTMOU�TT;RCVg? �SHELL_�WRK.$CUR�_STYL��Γ<OPT��?PT�B�?�2C�?R_DECSN_0<�L	O O-OVOQOcOuO�O�O �O�O�O�O�O_._)1�SSREL_ID�  ��Y�=UU�SE_PROG �%8:%*_�_>SC�CRk0ORY@3�W_HOST !8:#!�T�_�ZT\Ю_� c�_�Qc<o�[_�TIMEi2OV�U~)0GDEBUGMP�8;>SGINP_F�LMS`�gn�hTR\�o�gPGA�` �l�C�kCH�o�hTWYPE5<A)_ #_Y�}���� �����1�Z�U� g�y����������� ��	�2�-�?�Q�z�u� ������ϟ�
��eWORD ?	8;
 	PR�`�U�MAI@��3SU�1E�TE#`U���	�4R�COL�S�n���vTRACECTL 1��ŻB1 I�} ~�W d�ެ��_DT Q�����РD � *������W.��.��.���`.��"��	��
���
2�:�B�B����"���;���3�:�B� J��+�=�O�a�s���@������Ϳ߾��+Z��������#� ������������;� ��C���K���S���[� ����������,���Q��OP�����ą��\�nπ��� �Ħ ��������� � 2�D�V�h�zߌߞ߰� ���ߦ�q�3�E�W��� ��ϟϱ����_�� �%�7�I�[�m���� ������������! 3EWi��0\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz�u X����� �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� �ߚ������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�?��?OA�$PGT�RACELEN � A  ���@�$F_�UP ���e�SA[@?AT@�$A_CFG ��SE=CAT@��D�D�O�G6@�OhB�DEFSPD e�sLA6@�$@�H_CONFIG� �SE;C �@@dT�3B 	AQP�D�A1Q@ۂ$@INk@TROL �sM�A8�E�FQPE�E�W��SA�DQ�ILI�DlC�sM	�TGR�P 1�Yb@l�AC%  ��l��AA��;H�{N��R���A!P�D	� a3C	\�T�Ai)iQP� 	 �O4VGgCoG ´|c^oGkB` �a�opo�o�o�o�o�b"�Bz�o�7I~3 <}�<�oN�J� ����f�)��9�_�J�`z����@
t���d�ŏ�֏� ��3��W�B�{�f�x�@����՟�����J)@�)
V7.10�beta1�F �@�@ㅟA&ff�Q2�C�PC�`�D�Dk�`[�C�T��@ �DĠ Dr� ��QBH�`�L��PC�5R A?�  F��CCx����b��P`!P��A����Ap�By�b!PA1�������
�?L��?3�33A@��"��Fsff.��b�w:��7��AeC�QK�NOW_M  ��E{F�TSV �Z(R�C������ ʿ��ٿ�$�A!m�SM�S�[ ��B�	�E����Ϗ�̓E`��2�E@�2�������̭ L�MR�S�Y�T�j���AC5����e�@�Rۚ]ST�Q1 {1�SK
 4�U��A�¨߰E��*��� ��������J�)�;� M�_�q������� �����F�%�7�|��E�p�2{���A�<�����P3��������p�4��+p�A5HZl~p�6����p�7� $p�8ASewp�7MAD0F [Fp�OVLD  SK��ϼOr�PARNUM  /�O//_T_SCH� [E�
}'F!�)=C�%UP�DF/X)�/3Tp�_C�MP_O�0@T@@'�{E�$ER_CH�K5yH!6
?;RqS�]��Q_MO��o?�5_k?��_RES_GzФ~ݍ��? �OO�?%OO*O[ONO OrO�O�O�O�O�O�O��3���<�?_�5 ��(_G_L_�3G g_�_ �_�3� �_�_�_�3�  �_o	o�3@$oCoHo��3�co�o�o�2V �1�~կ1e�@c�?��2THR_ICNR�0�!7³5d�foMASS Zw�MN5sMON_�QUEUE ��~�f��0�� �4N�0UH1NEv6;�pE�ND�q�?�yEXE��u� BE�p��sOPTIO�w�;�p�PROGRAM %hz%�p�ol/~�rTASK_I���~OCFG ��h/\���DATA�Rè��@��2 �����#�5�G��k� }�������^�ן�������INFORé܍�wtȟe�w����� ����ѯ�����+� =�O�a�s���������hͿ(�4��܌ �Il��� K_�����T��ENB� ͻ1�>ƽ�I��G��2�~� P(O���ϳ� ������_EDIT ���ߋ�WERF�L�x�cm�RGADoJ �8�AС�i�?�0t�
qLֈq����5�?9�!��<@��*Ɓ%���@�#ߊ��2Y���F�	Hpl�G��b��>��A�d�t$I�*zX�/Z� **:c� �0V�h���Ǟ���B������������ ��������b���L� B�T���x��������� :����$,�P b������ �~(:h^p ������V/ / /@/6/H/�/l/~/�/ �/�/.?�/�/?? ? �?D?V?�?z?�?O�? �?�?�?�?rOO.O\O ROdO�O�O�O�O�O�O J_�O_4_*_<_�_`_ r_�_�_�_"o�_�_ooo�f	���o�p�o �o�dJ��oL��o#�o�GY��PREF S����p�p
L�?IORITY���}�P�MPDSP��>ߴwUTz�4�K�OoDUCTw�8��\�OG�_T�G;�|����rTOE�NT 1��� �(!AF_IN�E�pp�{�!t�cp{���!u�d��ˎ!ic�m�����rXY�Ӵv����q)� p�/�A��p�)�j�M� Y���}��������ן ���8�J�1�n�U�����*�s�Ӷ}}��毼��,�?:��jfBp�/z�֯K�,�������A��,  �p�������ʿ�u�"�ut�}�sF�P�PORT_NUM�s��p�P�_C?ARTREP�p�ξ|�SKSTA�w �K�LGSm���������pUn?othingϿ�������c{t�TEMPG ����ke���_a_seiban0C�,S�y�dߝ� ���߬�����	���� ?�*�c�N��r��� ���������)��M� 8�q�\�n��������� ������#I4m X�|�������3��VERS�I�p �d �disabled�>SAVE ���	2600H�721:&�!`;���̏� 	(H�rmoN+E/`�eb/ �/�/�/�/�*z,��? %`���_-� +1���E0�b�8eO?a?4gnpURGE_ENB3��v�u6�WF�0DO�v���vWi��4�q*�WR�UP_DELAY� �CΡ5R_HOT %�f�q:��.O�5R_NORM�ALH
�OrOAGS�EMIQOwO�OlqQ/SKIP-3���>3x$�O _1_C_] &ot_b_�_�_�_�_�_ �_�_o(o:o o^oLo �o�o�olo�o�o�o  $�oH6X~� �h��������D�2�h�z�����?$RBTIF�4G�RCVTMOU\������DCR�-3��I ��QE=o�C9�.E���C���A@_�8���J]ŦU�ŉ��mĚ�n´�?[����t_V�R_ ;��x5;��0;��i;�du;�t�<!��h��R���̝���� �&�8�J�\�n�����������RDIO_TYPE  4=���¯EFPOS1w 1�C�
 x/ :�H2��b�M���/�� E�οi�˿ϟ�(�ÿ L��pς��/�i��� ���ω�߭�6���3� l�ߐ�+ߴ�O����� �ߗ���2��V���z� ��9����o���� ���@�R�����9���������OS2 1��;+�u���-��xQ���3 1������G���gS4 1�~����ZE~�S5 1�%7q��/>�S6 1Ũ���/�/o/�/&/S7 1�=/O/a/�/?�?=?�/S8 1� �/�/�/0?�?�?�?P?�SMASK 1��߯ )�OF�7XN�OܯFUO_C�M�OTE���X4uA_?CFG �|M�1�\A�PL_RAN�GxA���AOWER� ���@�FS�M_DRYPRG %�%y?!_�ETART ��N�/ZUME_PRO��O_�_X4_EXE�C_ENB  <����GSPDdP�P8�X���VTDB�_�Z�RM�_�XIA_O�PTIONφ�����pAINGVERmS.a�z_��)I_AIRPU�R�@ @O�o�=MKT_�0T�@zO���OBOT_ISO�LC=N�F�1�a^�eNAMERl�bo��:OB_ORD_�NUM ?�H��aH721w  V1wLqrǈqrV0qr�sps�u\@��P?C_TIMĖ���x��S232�B1�����aLTE�ACH PENDcAN΀�7\H���x?c�Maint�enance C�onsV2�#�"��_�No Use��N��r�������8��С�rNPO>P�r�\A<e�qCH_�LgP�|Nw�	�<��!UD1:�b�	�R�0VAIL�Rq2e��upASRW  �:a�B��R_INTVAL1f��I�+n���V_DATA_GRP 2���qs0DҐP�?`��?�� o��������կï�� ���-�/�A�w�e� ���������ѿ�� �=�+�a�Oυ�sϕ� �ϩ��������'�� K�9�[߁�oߥߓ��� �����������G�5� k�Y��}������� �����1��U�C�e� g�y��������������	+Q?uDA��$SAF_DO_PULS�pE@�C��� CAN�r1f��vpSC�@�'��'Ƙ�Q�V0D��D�qL�L�+AV2  y�'9K]o��������ڈ���2($Md�($C!u�1#
) @�Co/�/�/�.W)k/� M��$�_ @݃T:`�/??�&?39T D�� 3?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO�jO|O֏��i%�O�O�O܉�!L� ��;�o݄�p��M
�t��D�ipp�L��J� � ��jL���j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:����/c�u������� ��Ϗ��B�%�1� C�U�g�y���������Ƒ��0RMS�EW] �$�6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ��M���*�<�N�`� r߄ߖߨ�������� ��&�8�J�\�ǟ�� �������������� ��,�>�P�b�p��� ������������ %7I[m�� �����!30EWit�OB3 t�����// //A/S/e/w/�/�/�/�/�/�*��/?6���\R?�M	�1234567�8XRh!B�!̺��� �?�?�?�?�?�?�? OOA�>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_o]-O�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�oq_BH�o�o�o !3EWi{���������v[;�j�A�S�e�w� ��������я������+�=�O�a�xYD� k�������ɟ۟��� �#�5�G�Y�k�}��� ����v_ׯ����� 1�C�U�g�y������� ��ӿ���	�ȯ-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� σߕߧ߹������� ��%�7�I�[�m������v6�����z��!�3�O:C�z  A�z  W �@�2�v0�� @�
���  	�r������X������ph�u�����K]o�� ������# 5GYk}��0 ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-?G��������*@  <X4t���$SCR_GRP� 1�'� �'�� t ��t� E5	 �1��2�2�4��W1G3�;�97�7�?�?OC���|�BD�` D���3NGK)�R-2000iC�/165F 56/7890��E��?RC65 �@�?
1234�E�6�t�A�����C �1F�1�3�1)�1A�:�1�I	��?_Q_�c_u_�_���#H��0 T�7�2�_��?�_�_o�6�t���_Lo�_poB8boK�h��@�UP{�  �$��1BǙ�B��  B�33BAƿ`�e�b�c�1Ag���o  @t��e�1@<>@	  ?�w�b�H�`2�j�1F@ F�`\rd[o� s������� *��9�a�a)rU�@�R�d�v�B����ʏ�� �ُ����H�3�l� W���{���Ě2C�?���7���9�t�:!q@"p>SԪD_��U�r�`y��`ȏ���G�L�3��ϯ�A >G�1��"oe��)	�t� �<�N�\��*�q�}���^� P��(����ӿ�g1�EL_DEFAU�LT  �D���t���HOTSTR� ���MIPOWERFL  K����?�oWFDO� S��RVENT 1�����P0� L�!DUM_EI�P翬��j!AF_INE��ϵO!FT������r�!�_B� ���i�!RPC_M'AINj�LغXߵ�N|�VIS��Kٻ����!TP��PU��߳�d��M�!
P�MON_PROX	YN��e<���g���f����!RD�M_SRV���g��1�!R�DM���Yh �}�!
~�M����il���!RL�SYN�@����8|��!ROS���<�4a!
C}E�MTCOMb���kP�!	vC'ONS���l���!vWASRCd ���m�E!v'USBF��n4� 0ߵ����/��'/�K//o/�RV�ICE_KL ?�%�� (%S?VCPRG1v/�*"�%2�/�/� 3�/�/"� 4??� 56?;?"� 6^?c?� 7�?�?�� \��?L19�?�; �$H�O�!�/+O�!�/ SO�! ?{O�!(?�O�! P?�O�!x?�O�!�?_ �!�?C_�!�?k_�!O �_�!AO�_�!iO�_�! �Oo�!�O3o�!�O[o �!	_�o�!1_�o�!Y_ �o�!�_�o�!�_{/�" � �/� F�E1�� ������
�C� U�@�y�d��������� �Џ����?�*�c� N���r��������̟ ��)��M�8�_��� n�����˯���گ� %��I�4�m�X���|������ǿ�ֿρ*_�DEV ����MC:�H~'�GRP 2ׇ��+p� bx 	_� 
 ,y�� ��+r~ϻϢ������� ���9� �]�o�Vߓ� z߷��߰������#� z�G���k�}�d��� ������������ U�<�y�`��������� *���	��-Qc J�n����� �;"_FX ��������/ �/I/0/m/T/�/�/ �/�/�/�/�/�/!?? E?W?�{?2?�?�?�? �?�?�?O�?/OOSO :OLO�OpO�O�O�O�O �O_^?�O=_�Oa_H_ �_�_~_�_�_�_�_�_ o�_9oKo2oooVo�o zo�o�o _�o�o�o# 
G.@}d�� ������1�� U�<�y����o��f�ӏ �̏	���-�?�&�c� J���n��������ȟ ����;���0�q�(� ��|���˯���֯� %��I�0�m��f������ǿ������R�d ��	�4��X�C�0|�gϠϯ�%�����R���������� �����+��O�=�s� ���Ϧ���i������� ���	��Q��x�� A����������� Y��P���)���q��� ��������1�U��� I��Ym��� 	�-�!E3 U{i���� ��//A///Q/w/ ��/�g/�/�/�/�/ ??=?/d?v?-?O? )?�?�?�?�?�?OW? <O{?OoO]OO�O�O �O�O�O/O_SO�OG_ 5_k_Y_{_}_�_�__ �_+_�_ooCo1ogo Uowo�_�_�oo�o�o �o	?-c�o� �oS�O���� �;�}b��+����� ����ɏ�ݏ�U�:� y��m�[�������� ş�-��Q�۟E�3� i�W���{����د� ��ï���A�/�e�S� ��˯���y��ѿ� ���=�+�aϣ���ǿ Qϻϩ���������� 9�{�`ߟ�)ߓ߁߷� ��������A�g�8�w� �k�Y��}����� ���=���1���A�g� U���y���������� 	��-=cQ� �����w��� )9_���O ����/�%/g L/^//7///�/�/ �/�/�/?/$?c/�/W? E?g?i?{?�?�?�?? �?;?�?/OOSOAOcO eOwO�O�?�OO�O_ �O+__O_=___�O�O �_�O�_�_�_o�_'o oKo�_ro�_;o�o7o �o�o�o�o�o#eoJ �o}k���� ��="�a�U�C� y�g�������ӏ��� 9�Ï-��Q�?�u�c� ��ۏ��ҟ������� )��M�;�q�����ן a�˯��ۯݯ�%�� I���p���9�����ǿ ��׿ٿ�!�c�Hχ� �{�iϟύ��ϱ��� )�O� �_���S�A�w� eߛ߉߿����%߯� ��)�O�=�s�a�� �߾��߇������� %�K�9�o������_� ����������!G ��n��7���� ��O4F� �g�����' /K�?/-/O/Q/c/ �/�/�/��/#/�/? ?;?)?K?M?_?�?�/ �?�/�?�?�?OO7O %OGO�?�?�O�?mO�O �O�O�O_�O3_uOZ_ �O#_�__�_�_�_�_ �_oM_2oq_�_eoSo �owo�o�o�o�o%o
 Io�o=+aO�s ���o�!��� 9�'�]�K�������� q���m�ۏ���5�#� Y�������I�����ß şן���1�s�X��� !���y���������ӯ 	�K�0�o���c�Q��� u��������7��G� �;�)�_�Mσ�qϧ� ���ϗ�ߓ��7� %�[�I���Ϧ���o� ���������3�!�W� ��~��G������� ����	�/�q�V���� ��w�����������7� .����O�s ����3�' 79K�o�� ����#//3/ 5/G/}/��/�m/�/ �/�/�/??/?�/�/ |?�/U?�?�?�?�?�? �?O]?BO�?OuOO �O�O�O�O�O�O5O_ YO�OM_;_q___�_�_ �_�__�_1_�_%oo Io7omo[o}o�o�_�o 	o�o�o�o!E3 i�o��Y{U� ����A��h�� 1�������������� �[�@��	�s�a��� ���������3��W� �K�9�o�]������� ����/�ɯ#��G� 5�k�Y���ѯ����� �{�����C�1�g� ����ͿW��ϯ����� ���	�?߁�fߥ�/� �߇߽߫�������� Y�>�}��q�_��� ������������ ��7�m�[�������� �������!3 iW������}� ��/e� ��U����/ �/m�d/�=/�/ �/�/�/�/�/?E/*? i/�/]?�/m?�?�?�? �?�??OA?�?5O#O YOGOiO�O}O�O�?�O O�O_�O1__U_C_ e_�_�O�_�O{_�_�_ 	o�_-ooQo�_xo�o Aoco=o�o�o�o�o )koP�o�q� �����C(�g �[�I��m������� ُ� �?�ɏ3�!�W� E�{�i�����؟� �����/��S�A�w� ����ݟg�ѯc��� ��+��O���v���?� ����Ϳ��ݿ��'� i�Nύ�ρ�oϥϓ� �Ϸ�����A�&�e��� Y�G�}�kߡߏ���� ���ߵ��߱��U�C�y�g����������$SERV_MA_IL  ������OUTPUT����RV �2؍�  � �(����_���SAV�E���TOP10� 2�9� d 	�������� +=Oas��� ����'9 K]o����� ���/#/5/G/Y/�k/}/�/�/�/���Y�P|���FZN_C�FG ڍ����j��!GR�P 2��'&� ?,B   A=0��D;� B>0��  B4��R�B21l�HELL��"܍�$�L�M��7�?�;%RSR �?�?�?O�?%OOIO 4OmOXOjO�O�O�O�O��O�O_!_3^�  �R3_a_s_AR_ ��{_�R�PS�xWIR2��d�\��]�Rh6HK 1�v; �_o"oo Fooojo|o�o�o�o�o �o�o�oGBT�fb<OMM ��v?�g2FTOV_�ENB��A�$��RO�W_REG_UI����IMIOFW�DL�pߥ~@5�WAIT�r�Y�8����v@�0�TIMn�u��j�VA��|A��_UNIT�s졆$�LC�pTRY��w$���MON�_ALIAS ?5e�yH�he��%� 7�I�[�i�������� m����
��.�ٟ R�d�v�����E���Я ������*�<�N�`� �q�������̿w�� ��&�8��\�nπ� �Ϥ�O���������� ��4�F�X�j�ߎߠ� �����߁�����0� B���f�x����Y� ����������>�P� b�t������������ ��(:L��p ����c��  �6HZl~) ������/ / 2/D/V//z/�/�/�/ [/�/�/�/
??�/@? R?d?v?�?3?�?�?�? �?�?�?O*O<ONO`O O�O�O�O�OeO�O�O __&_�OJ_\_n_�_ �_=_�_�_�_�_�_�_ "o4oFoXooio�o�o �o�ooo�o�o0 �oTfx��G� �����,�>�P� b����������Ώy�����(�:���$�SMON_DEF�PRO ����c� �*SYSTE�M*M�RECAL�L ?}c� (� �}7copy� frs:ord�erfil.da�t virt:\�tmpback\�=>192.16�8.56.1:7�360A�����}�.��mdb:*.*��ʞҟc�u����2x��:\,���>��0 V������3��a����T�ׯh�z� �������=�X���� � ���D�ֿg�yϋ� ��1�>�ԯ����	����Ͽ�R�c�u߇��
�xyzrate 61 .�@�R������������3700 ����d�v����0#�:picku�p.tp/�emp�=�<�T�����	��/��lace��0��� d�v�������6�I��� �����$Ͽ�����d v���,��<�V� �߯�>��h z���1CU���
/#�ϴ13924 ��e/w/�/�tpdisc 0-/? @/R/�/�/�?tpconn 0 �/�/�/a?s?�?8�����/?  �?�?�?�$�?7(�? dOvO�O,�:%WO�O�O_ 4#�O1. �Oi_{_�_�?�?;OVO �_�_oO�_BO�_eo wo�o�O/_A_�O�o�o _�o�oP_as�� 1�>P���1��4�4+�f� x�����,�?�X�U�� ��
�/��׀ď֏g� y����}.�@�R���� ��,���Пa�s��� �_�_3o�_߯��o (oïLo]�o����o�o ��oۿ���$�� 2�ڿk�}�Ϣ���=� X������ ���D����g�yߋߚ��$SN�PX_ASG 2���������  Y2%y�����  ?����PARAM ������ �	*��P������*�����OFT_K�B_CFG  ��ô՞�OPIN_�SIM  ���%������R�VQSTP_DS�Bk�%����SR� �� � }&��ONROD���0���TOP_O�N_ERR  �/�W�L�PTN ����A�H�RING_PR�MV� ��VCNT_GP 2��'��x 	������`�� ��$��VD��RP 1���(� ��_q��� ����%7 I[m����� ���/!/3/Z/W/ i/{/�/�/�/�/�/�/ �/ ??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_r_o_�_�_�_�_ �_�_�_�_o8o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c����� ������Ϗ���� )�P�M�_�q������� ��˟ݟ���%�7� I�[�m��������ܯ�ٯ����!�3�=P�RG_COUNT�L���[�_�EN�B��Z�M��N䑿_�UPD 1��T  
H���ۿ� ��(�#�5�G�p�k�}� �ϸϳ����� ���� �H�C�U�gߐߋߝ� ���������� ��-� ?�h�c�u����� ��������@�;�M� _��������������� ��%7`[m ������� 83EW�{� �����/// //X/S/e/w/�/�/�/ �/�/�/�/?0?+?=?�O?x?s?�?Q�_IN�FO 1�ɹ�� �F��?�?�?O�9��D�A���>>�O�3C+����BЁ@	��*7Ң¸�LY�T@P�YSDOEBUGi�ʰ�0�d��z@SP_PA�SSi�B?�KL�OG �ɵʴ��0>H�?  �����1UD1�:\�D�>�B_MPAC�Mɵ:_L_ɱ�A�j_ ɱVSAV ���MA�A�B�5� XSVnKTEM�_TIME 1��G�� 0��{r��rlXO  ���T1SVGUNS�İj�'���`A�SK_OPTIO�Ni�ɵ����?a_�DI�@��[eBC2_GRP 2�ɹ��T�o�1@�  C���cP��`CFG 3�k�\ b�k
}`
OB- Rxc����� ����>�)�b�M� ��q���������ˏ� �(��L�7�p����4m���n�ϟ�\��� ��;�&�_�q^�Qd T�������ѯ����� ��)�+�=�s�a��� ������߿Ϳ��� 9�'�]�Kρ�oϑϓ� �����Ȭ�����1� C���g�U�wߝߋ��� ���߳�	���-��Q� ?�a�c�u������ ������'�M�;�q� _��������������� 7��Oa� �!�����! 3EiW�{� ����/�/// S/A/w/e/�/�/�/�/ �/�/�/??)?+?=? s?a?�?M�?�?�?�? O�?'OO7O]OKO�O �O�OsO�O�O�O�O_ �O!_#_5_k_Y_�_}_ �_�_�_�_�_o�_1o oUoCoyogo�o�o�o �o�o�o�?!?Q c�o�u���� ���)��M�;�q� _�������ˏ���ݏ ��7�%�G�m�[��� �����ٟǟ���� 3�!�W�o������� ïA��կ����A� S�e�3���w�����ѿ ������+��O�=� s�aϗυϧ��ϻ��� ����9�'�I�K�]� �߁߷�m�������� #��G�5�W�}�k�� ������������1� �A�C�U���y����� ��������-Q ?uc����� ����/A_q ������/�� �$TBCS�G_GRP 2���� � �  
 ?�  J/\/F/�/ j/�/�/�/�/�/�/;�#"*#�1,d0�?1?!	 H�D 6s33�[2�\5O1B�x!x?�9D)�6�L�ͣ1>����g6�0CF�?�?�8fff�1�>��!OI/Cj��6�1H4?B�C{OO�)H��0|A�]0@HD�O_O)H�1�8CFr�O�M@ �. XU&_ �O_Q_n_9_K_�_�_��[?��0�Sp �	V3.00�R�	rc65�S	*`�T"o�V|A��0 8 `�Y �G`mHo  � ��%@�_�o�c#!J2�*#�1-�o�hCFoG ��;!�C!�j�B"]b�ox�BPz �Pva���� �����<�'�`� K���o�������ޏɏ ��&��J�5�n�Y� k�����ȟ������ \	��-�ן`�K�p� ��������ޯɯ�� &�8��\�G���k��� ��!/ۿ����� 5�#�Y�G�}�kϡϏ� ������������C� 1�S�U�gߝߋ��߯� ����	����?�-�c� Q���Y����m��� ���)��M�;�q�_� ���������������� %I[m9� ������! E3iW�{�� ���/�///?/ A/S/�/w/�/�/�/�/ �/�/?+?��C?U?g? ?�?�?�?�?�?�?�? OO9OKO]OoO-O�O �O�O�O�O�O�O_�O !_G_5_k_Y_�_}_�_ �_�_�_�_o�_1oo UoCoyogo�o�o�o�o �o�o�o	+-? uc����y?� ���;�)�_�M��� q�������ݏ���� �7�%�[�I������ ��o�ٟǟ����3� !�W�E�{�i������� ��ï�����A�/� e�S�u���������� ѿ�����+�a�� yϋϝ�G��ϻ���� ��'��K�9�o߁ߓ� ��c��߷�������#� 5�G���}�k��� �����������C� 1�g�U���y������� ����	��-Q? a�u����� ��/���q_ �������/ %/7/�/m/[/�// �/�/�/�/�/?�/? !?3?i?W?�?{?�?�? �?�?�?O�?/OOSO AOwOeO�O�O�O�O�O �O�O__=_+_M_s_ a_�_C�_�_}_�_ �_o9o'o]oKo�ooo �o�o�o�o�o�o�o #Yk}�I� �������� U�C�y�g��������� я����	�?�-�c� Q�s�u��������ϟ ��)�;��_S�e�w� !�����˯��ۯݯ� %��I�[�m��=������ǿ���վ  �� �)����$TBJOP_�GRP 2�ݵ��  K?��	A�H��O���� ����pX�d� ���� �� �,� �@�`�	 �D� ��Ca�D���`���f{ff��>��H����L��	�<!aM���>���=�?B�  Bp��8��C�D)�U�CQ�p�D�S�Ι㙚y���v� ?�������\<����U����%�C�V+��/���S�D5mi�{Բ��ع��<���z�>���\>�33C��  CA��`�K�j��u�bߐ���z��;�9bB��E�>�׵ҳ� C�V���s�����&��ǌ��;���6��%�]�D&� C��������
�>�� ?s33�����<Z;u���ff
�ҴK������U� )C-_i�u� �����*�IcM������Ƙ����	V3�.00f�rc65e�* e��/� ' F�  �F�� F� �F�  G� �GX G'� �G;� GR� �Gj` G�� �G�| G� �G�� G�8 �G�� G�< �H� H� �H��2 Ez  �E�@ E�� UEB F� FR FZ �F�� F� �F�P<"G � �GpL#?h G�V� GnH G��� G�� G��( =u=W+�(�$`QQ�?2�3�?�  ��M?[:A���*SYSTE�M
!V8.302�18 �38/1/�2017 A �y  p7M�T�P_THR_TA�BLE   $w $�1ENB��$DI_NO���$DO�4  ���1CFG_T � 0�0MAX�_IO_SCAN��2MIN�2_TI,�2DME\��0@��0  � �$COMMENT� $CVA�L	CT�0PT_I�DX��EBL�0N;UMQBENDIJfA�ZITID]B �$DUMMY13���$PS_OV�ERFLOW�u$�F�0FLA�0�YPE�2�BNC$?GLB_TM�7�E�F@�1�0ORQCT�RL�1�$DoEBUG�CRP�@�2@  $SB�R_PAM21_�VP T$SV�_ERR_MOD�U4SCL�@RAC�TIO�2�0GL_�VIEW�0 �4 $PA$Y*tRZtRWSPtR�A/$CA@A�1��_SUeU �0N|�P3@$GIF3@}$eQ lP_S�PNiQ LpP�VI<P��PF�RE�VNEA�RPLAN�A$�F	iDISTAN�Cb�1JOG_R�ADiQ@$J_OINTSP�ޤTMSETiQ � �WE�UACONqS2@B�RONFiQ�	� $MO�U1A`�$LOC�K_FOL�A�2B�GLV@CGL�hT?EST_XM@@ra'EMPE`,R�b�B`�$US;AfPH`�2P�S�a�bM�P_�`�aQCE�NEdRr $KA�RE�@M�3TPD�RAhP;t2aVEC�LE�32dIU�a�qHE�`TOOL�H`�0qsVI{sRE�SpIS32�y64N�3ACHX`�`~q3ONLE�D29�B�p�I�1  @$�RAIL_BOX�EHaPROBO��d?�QHOWW�AR�0�r�@�qRO�LM�B�A�C �SqK�r�@�0O_F9�C!��S�qiQ
>o� �RVpOCiQN_�SLOGaK��VKOUZbR�eA?ELECTE<P`��$PIP�fNOcDE�r�r�qIN�q�2^��pCORDE!D�`�`}��0P9P@  D �@OBAU`TA�a� ���C�@���P�q0���ADRA�0F@TC}Hup  ,�0SEN�2�1A�a_�T�l�Z@�B�RVWV�A!A � �ApeR�5PREV_�RT�1$EDI}T��VSHWR9��S@	UАIS`yQ/$IND0@1QB�~�q$HEAD�`5@ ��p5@��KEyQ��@CPSPD�J�MP�L�5�0RA[CE�4�a��It0S�CHAN�NEzp�	WTIC�K{s�1M`A�0@�H-N�AD0^�]D��`CG�P���v�0S3TYf��qLO�A�3�B���jP t 
���Gr�%$���T=�PS�!$UN�IGa5A�E�0�FPO;RT��SQU5ptR��B�TERC�J@���TSG�� �PP6�$�DE$��$`Thq�0OK@>CFV�IZ�D�Q�E�A�PR�AͲ�1��P9U}aݵ_DObk��XSV`K�6AXIt��7�qUR_s��E$T�p��*��0F�REQ_hp<�ET�=�P�b�PARA�`@.P
@�[���ATHr�3@�D�s�sv�0 �2SR_Q��0l}��@�1T�RQIc��$`�@��B�Rup��VE@@��NOLD��Ap7a���x@�A��AV_M�G�����/���/�D�)�D;�DM�J_AKCC.�C��<�CM��0CYCM@3@��M@�_E�����٘@�NbSSC�@  hPDS���1�@3SP�0*�AT:�����@��i��BADDR�ES{sB��SHIyF}b�a_2CH�@�&�I�@|��TV
�bI�2]��h>��C*�
�j
�2V���N�0 \��������웱�@��CnӞ�a��ꯆ:R���TXS�CREE��0�TINAWS�P;�ºT�1>�>�jP TQ�7P�B�6QP���
��
���RROR_"a�@���D�1;UEG� ���U�r�@SXQ�RSM�� �UNEXg��6���0S_�S��	�0��>�C�b��o� �26�UE����2GRUͰGMT/N_FLQ�#P�OHgBBL_�pW�g@�0 ����O�Q�LEn���p�TO`C�RIGH��BRDITd�CKsGRg@�TEX,�|��WIDTH�s�ݐB�A�A{q��I�_/@H��  o8 $LT_ �|�Y0@RyP�b�s�wH�B��GOu��0D0ITW� U� �R�b��LUM�!�^�E#RV��]PFP`>���1'@r�GEU�R�cF\��Q)��LIP�Z�Ed��)'@�$(�$(�p#)5!+6!+7!+8"b�>C�Ȱ`��F�q�aSv�@EUSReTO  <��/@U�R���RFOChq�PP�RIz�m�@?A� T�RIP�qm�U)N�0�4!�P ��0��5�7��b;�5� q"T� ̱G �aT7���}�O2OSNA�d6RA���;3wq�1#�n_�S�^�2�����aU!"A$�?�?+"��N;3OFF�` P%O���3O@ 1#�PD,D$PGUN�#K`S�B_SUqBBPk SRT�0�&��"avp��OR��p�ERAU���DT<�Ib��VCC��H��' ��C36M�FB1��PPG�?�( (b`�STE�Qʀ9PWTѠ�PE���GXd) y����JMOVE��{Q6RAN4`?[�3DV|�S6RLIM_X�3 qV�3qV\XvQk\:V01�IP�2VF��C!砽@��G�*���IB�P,�S� _��`�p�b���@ (0GB�� "P�@��|pr+x �r �,�tRn@��s 9C@TeDRI�PSfBQV!�wdԐ��D�$?MY_UBY�$\d �;QA�S���h�q��bP_S�ף�bL��BMkQ$j�DEYg�EX� ���B_UM_MU6�X�D<q US�?��;V=Go�PACI�TP �<Uyr�3yrkSyr:�;qREnr�1l��9cyr�@,�BTARGPP�p�R<a9R{0�@- d���;cB	:r��R�DS�Wqp�Sn�:s˰OD�!d�Av�3���E���U�p0m��vHK
�.��K�AQ��0�̍�?SEA����WO�R�@3��uMRCV�r/ ��O��M
�@C�	ÂC�sÂREF��̆��gR j�
�� Ȋ�ي��8=�̆r�_RC��s� ����@����b����sY�to0 �Т��;��� �e�OAU���r��\c(`+�u���2��<���̰� �-=���f�K�SU�L3a.�C7Po/+p�NT�a��]���ag��g��!g�&�L��c���c������!R�@T��s�1���>o@AP_HUR�ۥ�SA>SCMP��FP�����_&�R�T�������X.���V�GFS�E2d ��M� � Y0UF�_�����J��RO`� ����W,rUR�#GR�mq�I���D_V_h[D�@zY��3�WIN.rH���X-�V
A�RqR�P�W Ew�w�q|c6v,q��RvLOiPtc�PMc���3t +=�PA�' =�CACH 6����ŵ�,p��2K�jۓC�QIo�FR"�qT� $֭�$HO�@�R��`�rc��[�`֘p��ڔ�VP�r<����_SZ3p���6����12� ��]pآ؆P��WA3�MP\��aIMGx����AD�qIMRE�ٔ6�_SIZ�P���!po�6vASYN�BUF6vVRTD�h�t�F�OLE_C2D�T��t��0C0a�Us��QP�X�EC;CU�xVEM�p��<��#�VIRC��VTP�����G�p���t��LA�s�!����Mco4��;�C/KLASQC	��ђ�@5  �A�� �@&B�T$��$`��6� |F@o���Xñ�T@�o�?a��"�uI��جr/��`BG� VEJ�`PK|p1���֖�K�MHO+��R7 � }F���E�SLOW}w]RO>SACCE*@-�=�xVR:��11�yrcAD�/0rPA�ԩ&�D�1�M_qBa�81��JMP����A8y�b�$SS�C6u��M��C��@9$2��S8��N/�PwLEX��: T��C�Q��6�FLD6?1DEZ�FIQ r�O�qty� K�P}2��;� ϱ�PV多�MV_PIZ��G�BP��`а&�FIQ�PZ�$��������G9A%p�LOO0Tp�JCBT*����� ��ړPLAN�R&�L�F���cDV�'AM�p���U�$�S�P .q�%�!�%#�㱶C�4G����RKE<�1�VANC]K�\A0p <�@�?��?Q3A�a =��?q??T0�9��r># hܰ�	��K9�fdA2b<X@̠OUe��ݒA��
O���SK�(�M�VIE�p2�= S0:�|R?� <{@X���`UMKMY����Re��mD��ȧCU�`zb�U�@@ $�@�TIT 1$P�R8�UOPT��VSHIFʀ�A`�a���D�0�����$�_R$�U ړQ.qZ�U�s�o@t�Qav�Q5fSTG@�cVSCO��vQCNT���3� }w�RlW�R zV�R�W�R�XLo^opj*jA2��51D>a�0�� �pSMO"��B%TC�J�@1uK���_���@C%�Gi�LI� '�/�XVR�DDY�@�T��ZABCP�E�r�b���]
�ZIP�EF%���LV��L���^�bMPCF�eGy��$p	�rDMY_LN$@Ar8��dH ���g��>��MCMİC��CA�RT_Xq�P�1 �$JvsptD ��|r�r�w���u����UXW�puUXE#UL�x�q�u�t�u@�q�q�y�q�vJ�Z�eI Hk�d����Y�`D�� J �8o�	V�EIGH���H?("��f��ĔK �= �C����`$B&�K���1_X�B��LgRV� F�`��COVC؀qrfq 9��@}�e�
�����7�D�TRȰ	�V��1�SPH� ǑLa !�S�i�{�����ST�S  g��������a v�<�ѐNa1 ��w�� ����������������������"��	���a������
����������( N��RDI������@ğ֟����t�O|����������ίஔ�Sz��� >�����ſ׿ �����1�C�U�g� yϋϝϯ��������� �v�}���8�!�3�E� W���'�9�K�]���l� ����U��� ��( ��N� ��@A�|v�^`BF_TT��ի���I�V>0n�J�z_�I�R 1&� 8����%к� ��C�  ����� �������"�4�F�X� j�|������������� 1gBTjx�����р�����0B QI �ZlJ����� ����/"/4/F/ X/FҒ�t/�/b*���/P�/��bv�@`�v�MI_CHANU�E `� #3�dV�`�쓑&0ET>�AD �?��y0�m�@�/�/�?�?�d0RLP6s�!&�!�4�?~�<SNMASKn8|��1255.4E�0�33OEOWO�OO�LOFS^Q  ��%X9ORQCTROL &�V�m��O��T�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo(l�OKo�:ooo��PE�pTA�IL8�JPGL_C�ONFIG 	��ᄀ/ce�ll/$CID$/grp1so�o�o1�#��?\n ����E��� �"�4��X�j�|��� ����A�S������ 0�B�яf�x������� ��O������,�>� ͟ߟt���������ίB�}c���(�:�L� ^���`o��e��b��� Ϳ߿���\�9�K� ]�oρϓ�"Ϸ����� �����#߲�G�Y�k� }ߏߡ�0��������� ���C�U�g�y�� ���>�������	�� -���Q�c�u������� :�������); ��_q����H ��%7�[�m����]`��User V�iew �i}}1�234567890�
//./@/R/Z$X� �cz/���2� W�/�/�/�/??u/�/�3�/d?v?�?�? �?�??�?�.4S?O *O<ONO`OrO�?�O�.5O�O�O�O__&_�OG_�.6�O�_�_�_@�_�_�_9_�_�.7o_ 4oFoXojo|o�o�_�o�.8#o�o�o0�B�ocir l�Camera ��o������NE�,�>�P��j��|�������ď�I   �v�)��&�8�J�\� n���������ڟ� ���"�4�[��vR9 ˟��������ȯگ�� ���"�m�F�X�j�|� ����G�Y�I7���� �"�4�F��j�|ώ� ٿ����������߳� Y�����Z�l�~ߐߢ� ��[�������G� �2� D�V�h�z�!߃unY� ������������B� T�f������������ ����Y�"i{�0BT fx�1���� �,>P��Y� �i������� �/,/>/�b/t/�/ �/�/�/cu9H/�/ ?!?3?E?W?�h?�? �?F/�?�?�?�?OO/O�j	�u0�?jO|O �O�O�O�Ok?�O�O_ �?0_B_T_f_x_�_1O CO�p�{._�_�_oo +o=o�Oaoso�o�_�o �o�o�o�o�_�u�� �oOas���Po ���<�'�9�K� ]�o�PEc����͏ ߏ����9�K�]� ����������ɟ۟�� ��ϻr�'�9�K�]�o� ��(�����ɯ���� �#�5�G��;�ޯ ������ɿۿ��� #�5π�Y�k�}Ϗϡ� ��Z�����J����#� 5�G�Y� �}ߏߡ��π������������  ��N�`�r�� ������������   $�,�J�\� n��������������� ��"4FXj| ������� 0BTfx�� �����//,/�>/P/b/t/�/�  }
��(  �B�( 	 �/�/�/ �/�/??8?&?H?J?�\?�?�?�?�?�?�*4� �n�O1OCO ��gOyO�O�O�O�O�� O�O�O_VO3_E_W_ i_{_�_�O�_�_�__ �_oo/oAoSo�_wo �o�o�_�o�o�o�o `oroOas�o� �����8�'� 9��]�o��������� �ۏ���F�#�5�G� Y�k�}�ď֏��şן �����1�C�U��� y��������ӯ��� 	��b�?�Q�c����� ������Ͽ�(�:�� )�;ς�_�qσϕϧ� �� ������H�%�7� I�[�m���ϣߵ��� ������!�3�E�� ��{����������� ����d�A�S�e��� ������������*� +r�Oas��8����0@ �������� ���)frh:\tp�gl\robot�s\r2000i�c6_165f.xml�`r��������/����/3/E/W/i/{/�/ �/�/�/�/�/�//
? /?A?S?e?w?�?�?�? �?�?�?�??O+O=O OOaOsO�O�O�O�O�O �O�OO_'_9_K_]_ o_�_�_�_�_�_�_�_ _�_#o5oGoYoko}o �o�o�o�o�o�o o�o 1CUgy�� �����o��-� ?�Q�c�u����������Ϗ��K �� 88�?��2��.�P�R� d����������П� ��(�R�<�^���r������ܫ�$TPG�L_OUTPUT� ���� ����%�7� I�[�m��������ǿ ٿ����!�3�E�Wπi�{ύϟϱ������ˠ2345678901�������� 0�8�����_�q߃ߕ� �߹�Q߽�����%�7���}A�i�{��� ��I�[�������/� A���O�w��������� W�����+=�� ��s�����e �'9K�Y �����as� /#/5/G/Y/�g/�/ �/�/�/�/o/�/?? 1?C?U?�/�/�?�?�? �?�?�?}?�?O-O?O QOcO�?qO�O�O�O�O�OyO֡}�_)_;_M___q_�]@��_�_�� ( 	  ���_�_o�_5o#oYo Goioko}o�o�o�o�o �o�o/UCy g��������	�?��Ƭ�-�G� u���c�������ߏ� ��`��,�ΏP�b�@� �������Οp�ޟ� ���:�L���p���$� ������ܯ�X���$� Ư�Z�l�J������ ƿؿz�����2�D� ��0�zό�.ϰ��Ϡ� ����b��.���R�d� B�tߚ������߄� ����<�N��r�� &��������Z�l� &�8���\�n�L����� �����|�����  FX��|�0�� ���d0�  fxV���� �//�>/P/�</ �/�/:/�/�/�/�/?�
2�$TPOFF_LIM [��@W����A2Nw_SV#0  �T�5:P_MON �S�74�@�@2�U1STRT?CHK S�56�_=2VTCOM�PATJ8�196VW�VAR j=\�8N4 �? O�@}21_DE�FPROG %��:%CONRO�D�6kO�6_DIS�PLAY*0�>?BI�NST_MSK � �L {JIN�USER�?�DLC�K�L�KQUICK�MEN�O�DSCR�EPS��2tpsc�D�A1P6Y452GP_KYST�:59�RACE_CFGS �Fr1�4.0�	D
?��XHN/L 2�93��Q�; $B�_�_o o2o�DoVohozj�UITE�M 2�[ ��%$123456�7890�o�e  �=<�o�o�os  #!{!@�oZ C�o{�o��� 9K�o/��?�e� �����#���G� ��+���O���ŏ׏ Q�����͟ߟC��g� y����]��������� ���-���Q��u�5� G���]�ϯ!����ſ )�տ���q�ϕ��� ��3�ݿ�ϯ���%��� I�[�m���	ߣ�c�u� �ρ������3���W� �)��?���ߌ��� ������c�S�e�w� ������k������ ��+�=�O���s�E W��c������ 9�o��n �����#�G �"/}=/�M/s/�/ ��///1/�/U/? '?9?�/]?�/�/�/i? �??�?�?Q?�?u?�? PO�?kO�?�O�OO�OP)O;O_�TS�R�_>UJ�  �bUJ� �Q`_UI
 �m_�_z_�_8ZUD�1:\�\��QR_GRP 1�k�� 	 @ `@o!koAo/oeoSo�own��`�o�j�a�_��o�o�e?�   '9{#YG}k� ���������C�1�g�U�w���	��E��ÏSSCB ;2%[ � !�3�E�W�i�{������\V_CONFIG %]�Q]_�_����OUTPUT� %Y�����S�e�w������� ��ѯ�����+�_A @�S�e�w��������� ѿ�����+�<�O� a�sυϗϩϻ����� ����'�8�K�]�o� �ߓߥ߷��������� �#�5�F�Y�k�}�� ������������� 1�B�U�g�y������� ��������	->� Qcu����� ��);L_ q������� //%/7/H[/m// �/�/�/�/�/�/�/? !?3?D/W?i?{?�?�? �?�?�?�?�?OO/O AOݟ�>�O�O�O�O �O�O�O�O_!_3_E_ W_J?{_�_�_�_�_�_ �_�_oo/oAoSod_ wo�o�o�o�o�o�o�o +=Oaro� �������� '�9�K�]�n������ ��ɏۏ����#�5� G�Y�j�}�������ş ן�����1�C�U� g�x���������ӯ� ��	��-�?�Q�c�t� ��������Ͽ��� �)�;�M�_�p��ϕ� �Ϲ���������%� 7�I�[�m�~ϑߣߵ� ���������!�3�E��W�i�LH��� ����s���hO���� ��1�C�U�g�y��� ������t�����	 -?Qcu��� �����); M_q����� ��//%/7/I/[/ m//�/�/�/�/��/ �/?!?3?E?W?i?{? �?�?�?�?�?�/�?O O/OAOSOeOwO�O�O �O�O�O�?�O__+_ =_O_a_s_�_�_�_�_ �_�O�_oo'o9oKo ]ooo�o�o�o�o�o�o �_�o#5GYk }������o� ��1�C�U�g�y����������ӏ���$T�X_SCREEN� 1�����}��&�8�J�\�n������� ��ҟ��������� P�b�t�������!�ί E����(�:�L�ï p�篔�����ʿܿ� e�w�$�6�H�Z�l�~� ��������������  ߗ�D߻�h�zߌߞ� ����9�K���
��.� @�R���v��ߚ����������k���$U�ALRM_MSG� ?���  ��zJ�\��������� ����������/"S�Fw+�SEV  ��E��)�EC�FG ���  �u@� � A�   B��t
 x�s� 0BTfx������GRP �2� 0�v	� �/+�I_B�BL_NOTE ��
T�G�l�r��q� ~+"DEFPRO5�=%9� (%k�/ �p�/�/�/�/�/?�/ %??6?[?F??j?�?�!,INUSER � o-/�?I_M�ENHIST 1|8��  (| � ��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1�?`OrŌO�O�)'O9N381,23�O�O�O	_�O+�O9Eedit~EBCONRODMO�i_{_�__&O�O138,2�_�_�_o"o<�_�_,166X_no�o�o�o�@-7oA_SR2,1^o�o
'o�o;N4]ov����@'?Q~2LO�
� �.�Q#�0"A�?_�q� ���������CN���� ��+�=�̏a�s��� ������J�ߟ��� '�9�ȟڟo������� ��ɯX�����#�5� G�֯k�}�������ſ T�f�����1�C�U� @�yϋϝϯ������� �	��-�?�Q�c��� �ߙ߽߫�����p�� �)�;�M�_�q� �� ���������~��%� 7�I�[�m�������� ����������!3E Wi{fϟ��� ��/ASe w������ /�+/=/O/a/s/�/ �/&/�/�/�/�/?? �/9?K?]?o?�?�?"? �?�?�?�?�?O#O�? GOYOkO}O�O�O�:O �O�O�O__1_4OU_ g_y_�_�_�_>_�_�_ �_	oo-o�_�_couo �o�o�o�oLo�o�o );�o_q�� ��HZ���%� 7�I��m���������Ǐ�J�$UI_P�ANEDATA �1������  	��}/frh/c�gtp/whol�edev.stm�ӏ1�C�U�g�R�)Gpri���]�}���Ɵ؟���� � ) "�F�-�j�Q������� į��������B��T�;�x�V����     rP����ǿٿ ����b�3Ϧ�W�i� {ύϟϱ�������� ���/�A�(�e�L߉� �߂߿ߦ���������� ��8���T�Y�k� }�������J��� ��1�C�U���y��� r�����������	�� -QcJ�n� �0�B��); M�q����� ��/h%//I/0/ m//f/�/�/�/�/�/ �/�/!?3??W?�� �?�?�?�?�?�?:?O O�AOSOeOwO�O�O O�O�O�O�O�O_ _ =_O_6_s_Z_�_�_�_ �_�_�_d?v?4O9oKo ]ooo�o�o�_�o*O�o �o�o#5�oYk R�v����� ��1�C�*�g�N��� ��o"oӏ���	�� -���Q��ou������� ��ϟ�H���)�� M�_�F���j������� ݯį����7����� m��������ǿ�� ��p�!�3�E�W�i�{� ⿟φ����ϼ����� �/��S�:�w߉�p�`�ߔ���D�V�}���@�-�?�Q�c�u�)	� ��ŉ����������  ���D�+�h�O�a��� �������������@R9v	�`�Z���$UI_POST�YPE  `��� 	 ����QUICK�MEN  ����� RESTO�RE 1 `��  ��i�S`N�m ~������/ %/7/I/[/�/�/�/ �/�/r�/�/�/j/3? E?W?i?{??�?�?�? �?�?�?�?O/OAOSO eO?rO�O�OO�O�O �O__�O=_O_a_s_ �_(_�_�_�_�_�_�O �_o"o�_Fooo�o�o �o�oZo�o�o�o# �oGYk}�:o� ��2���1�C� �g�y���������d�����	��-��SC�RE� ?��u1scHuU2h�3h�4h�5h��6h�7h�8h��UGSERJ�O�a�TI��j�ksr�є4є5*є6є7є8ё� �NDO_CFG �!����Ѩ PD�ATE ����None _�� ��_INFO �1"`�]�0% 3�x�	�f�����˯ݯ ������7��[�m��P�������ǿ�J�O�FFSET %�ԿσA֏�*� <�N�{�rτϱϨϺ� Ͼ����A�8�J߀w�n߀ߒ�����
�����UFRAM/E  ʄ�G��RTOL_ABRqT&��>�ENBG�~8�GRP 1&<�Cz  A� ������������ ����:�� Ug��~V�MSK  j�]�X�N#���]�%x�߫��VCCM��'���RG��*��	��ʄƉD. � BH)�p<2�C�)��PN?�l` ��MR��20��Pp���"�р	 ����~XC56 *Ȩ�����N�5�р�A@<C�N ��� ʈ);h�c��Rр|�Ђ B���� 6�t/T1/ /U/ @/y/d/�/�/�/�/*/ �/	?�/???�c?u?.��TCC��1��f��9�рр��G�FS�22w �Й�2345678901�?�2ʈ"� 6��?!Oс>,12�QO�_GB@R 8N:�o=L��� ��������OOA �O�O@O_dOvO�O�O �O�_�O�O�___�_ <_N_`_r_Soeo�_Ro �o�_�_oo&o8o�>�4SELECF�j��$�VIRToSYNC� ���6�BqSIONTM�OU-tр���cu��3U��U��(�� F�R:\es\+�A\��o �� M�C�vLOG�  � UD1�vEX��с' B@� ����q  �ESKTOP-8U37T7F�6�!��N�`��3�  =�	 1- n?6  -��ʆ��xf,p�#�0=�̩ʹ���r�xTRAIN��2�1.���
. d��sq4w (,1��0�� )�;�M�_�q������� ��˟ݟ���I���crSTAT 5���� ������'$���ۯ�_GE��6nw�`. �
���. 2�HOMIN���7U��UC� �r�a�a�aCG��um�JMPER�R 28w
  �oE:��suTs���� �߿���'�9�OϠ]ώρϓ�_v_�pR�E��9t���LEXr��:wA1-e��VMPHASE � RuCCb��OcFFLpc�<vP2�t�;4�04��8����b@��ab>?Gs33��Á�1�рL��ҕԈ�|��t�>�x��Â��C{A�SDE�R-���o��E�B���-
.?O�W�  �E�4�B�� 2ҠƘ��� �^���0��<�1�`� ��� `�r�������>���� L�>��Jtn ������ �$6 �&4F\��� ����j// 0/Z/��\/��/�/ ��/T/�/ ??d/Y? �/z?�/�?�/�/,?�? �?�?ON?COr?�?�? �O�?`OO�O�O�O_ 8O�O_nOc_u_�O�_  _�_�_�__o4_&o X_Mo|_�_�_~o�o�o��o�g��TD_FI�LTEt�?�� ��Wp��]o$6 HZl~���� ����)�;�M��_�q������SHI�FTMENU 1-@x�<��%��� ��я��0���f�=� O���s�����䟻�͟����P�'�	L�IVE/SNAP�D�vsfliv��b���IO�N G�U���menu����:������l����A���	����b�K��5M���)�@�����A�pB8������Ӝѝ�r�����m`� ;�,��/�ME��u��Y�᱁MO��B����z��WAITD_INEND�3����OKN�.�OU�T#��Sa�4�TI]M�����G� ��@���`ϱ�ϱʞ��2�RELEASE�����TM���=��_ACTx������2�_DATA C�ի�%i��ߪ����RDIS�b�_�$XVR2�D���$ZABC_G_RP 1E8�n`�,@h2��ǽZIP1�FD� cCo�������x�MPCF_G 1G8�n`0<o ����=�H8����t� �	�w�  8�R�����e�����?� k������5��
\���  � a �����7������I��z��YL�IND�aJ�� ��f ,(  *s�K�p���� �//+.m N/�r/Y/k/�/��/ �/�/3/?�/�/J?1?�n?U?�/�?�?v�C�29K8��� ��O `o�7O~[Ol�?�O�g��AA�ASPHERE 2LS�?�OX?�O__>_ �?�Ot_�_?�_I_/_ �_�_o�_]_:oLo�_ �_�o�_�o�o�o�o#o� $7�ZZ� �k�