��   ��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_�$$C�LASS  ������D��D�VERSION�  ��
/IRTUA�L-9LOOR� G��DD8�?�������k,  1 <DwH8G�����D'�82 ��-��Z�Z]/o/�/ S/�/�/�-_ �/�/|�/;�$MNU>)AP"�� 8�'/ �!I?�?m??�?�? �?�?O�?O7O!OCO mOWOyO�O�O�O�O�O��O_�'5NUM � ��>�\P<UT�OOL/?4 
�E;U�P���.bQ3�P�Q��C�_ #_�_�O�_o�_o7o !oComoWoyo�o�o�o �o�o�o�o�o-W�Ac�9XiQIVyWV�