��   ��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_  �$$C�LASS  ������D��D�VERSION�  ��
/IRTUA�L-9LOOR� G��DD8�?�������k,  1 <DwH8G�����D'�82 ��-��Z�Z]/o/�/ S/�/�/�-_ �/�/|�/;�$MNU>�AP"�� 8����͋����T=P0K13���}2�o������)!D�_�?��C� #� �?�?�?�?�?�?O �?O7O!OCOmOWOyO �O�O�O�O�O�O_�~'5NUM  ���>�w%2TOOL�/?4 
E4,�^P���.Q3�P�Q��C�_#_�_�O �_o�_o7o!oComo Woyo�o�o�o�o�o�o �o�o-WAc��9XiQIVyWW�