��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�   � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d PPINFwOEQ/ ��L A �!�%/� H� �&�)EQUIP 2� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CE�S0s!_81s!9�K2> �! � �$SOFT�T�_IDk2TOTAoL_EQs $�0�0NO�2U SPI�_INDE]�5X�k2SCREEN_�(4_2SIGE0�_?q;�0PK_F�I� 	$TH{KYGPANE�4� � DUMMYE1dDDd!OE4LA�!R�!R�	 � $TIT�!$I��N �Dd�DPd �Dc@�D5�F6�FU7�F8�F9�G0�G��GJA�E�GbA�E�G1P�G �F�G1�G2�B~!SBN_CF>"�
 8F CNV_�J� ; �"�!_CM�NT�$FLA�GS]�CHEC��8 � ELLSE�TUP � 7$HO30IO�0� �%�SMACRO��RREPR�X� D�+�0��R{�T UTOBACKU��0 �)DoEVIC�CTI*0��� �0�#�`B��S$INTERV�ALO#ISP_UsNI�O`_DO>f<7uiFR_F�0AIN�1���1c��C_WAkda�jO�FF_O0N�DEL�hL� ?aA�a1b�?9a�`C?���P�1E��#sATyB�d��MO� ��cE D [Mp�c��^qREV�gBILrw!XI� ~QrR  � �OD�P�q$NO^PM�Wp�t�r/"�w� �u�q�r�0D`S p{ E RD_E�p~Cq$FSSBn&�$CHKBD_S�E^eAG G�"?$SLOT_��2$=�� V�d�%��3� a_EDIm  ? � �"���PS�`(4%$EyP�1�1$OP�0r�2�a�p_OK�;UST1P_C� ���d��U �PLACI�4!�Q�4�( raC�OMM� ,0$D ����0�`��EOWBn�IGALLOW�G (K�"(2�0VARa��@�2ao��L�0OUy� ,�Kvay��PS�`�0M�_O]����C�F�t X� GR�P0��M=qNFL�I�ܓ�0UIRE��$g"� SWIT{CHړAX_N�P]Ss"CF_�G�� �� WARN�M�`#!�!�qPLI��I�NST� CO�R-0bFLTR^C�TRAT�PTE�>� $ACC1a��N ��r$ORIأo"��RT�P_S�Fg CHG�0I���rTא�1�I���T�I1��� x i#�Q��HDRBJ; C,�U2'�3'�4'�5'�U6'�7'�8'�9s!uӡO`T <F �П����#92��LL�ECy�"MULTI�b�"N��1�!����0T_}R  4F STY�"�R`�=l�)2`�����`T |� �&$c��Z`�pb��P�MOL�0�TTOӰ�Ew�EXT����ÁB����"2� ��[0]�}R���b�}� D"}��� �Q���Q�kcG��A�^ȇ1��ÂM���P�� ŋ� L�  ���P�z�`A��$JOBn�x/�i�G�TRIG�  d�p�߻��� ��7��������_�M�b! t�pF̝ CNG AiBA � ����M���!���p � �q��0��P[`��,i�*�"6���0t�B񉠎"J��_Rz�gC�J��$�?�Jk�D�%C_�;������0ФR�t#�C ������G����0NHANC̳$LGa��B^a��� �D��A�`��gzRɡ�!��p�3DB�RA�sAZ�0KELT��\���PFCT&��1F�0�P��SM��cI��1�% ��% ��@R��a���� S��&���M 00{o Ve#HK~�A^S��h�����I_T$�"�6SW�CSXC�)�?!%��p)3��T�$@��PANN�&�AIMG_HE�IGHCr�WIDLI AVT�0��H F_ASPװ��`�EXP�1���CWUST�U��&��
|E\�%�C1NV q_�`�a��' \%1y�`OR�c,"�0gsdk��PO��LBSYI�G��aR%�`좔Psp�m��0k�DBPXW�ORK��(��$�SKP_�`ma1D�B<qTRp ) ���P���� �0f�DJ!d/�_CN�0�R�#� �'PL�S�Q��d�s�DKA7WA w'�^A�@NFZpfB�DBU��*�"!P	RS�7�
ЖQ����g+ [pr�$1�$ZϢ�Li9,�v?�3ʠ��-�?�4Cr��.�?�4ENEy���� /�?�3J0R�E`��20H��C�uR+$L,C,$pi3
�? =KINE@�fK!_D�I�RO�` ����ȳqvC��h ��FPAÃ3uR�PRYN�B�MR��U!�vu�CR[@EWM ^�SIGN��A�� .q�E�Q-$P���.$Pp 2�	/ P7�PT2�PDu`L���VDBAR@�GO_AW���Jp� ��DC�S�pZ�CY_ �1���@1<�Q?fI+G2�Z2>fN>������
�qS&c}P2 P7 $��RB?�e�eP=hPwg�QBYl��`gT+1�THNDEG�23��KS�SE|�Q��SBL�Y�ccҙT�!sQL�4� HpZ ���VTO3FB�l�FEfA��пb�TqSW5�bDO8C���MCS�f�`PZ$r�b H� W0�z�T�eSLAV�1;6�rINP��f���LyqQP�7� $,�S���=��vX��uFI��r@줭sc�!��!W1�N�rNTV'��rV	�n�uSKIvTE�@`W���:�J_�� _�00�SAFEܡA�_SV��EX�CLU��B �PDJ L1�k�Y�d�ƻ�rI_V� !PPcLY 0b���DE~wΙ�_ML2�B $�VRFY_�#��Mk�IOU��憻 0�d��:�O�P��LS�@�jb;�3572��Sr�� Px%X�{P�hs�� �� 8 @� T�A� qঠ ^�c_SGN��96� ���@�A�����iP`t!��s"��~UN�0@jdՔ�U���B �@ � ��� ���g��W I�2: @�`Fؒ���OT�@@�:4H1(�774C2�M`NI�2;�R�������A�q��DAY1#LOAD�T/4~�;30�o �EF�XI�b%< @%1O㠈3�� _RTRQ��=� D�`@��Q@  �EjP"�㥎��<�B�� 	�@��A#MP��]>�a�`����a�8Sq�DU�@�q���"CAB��?�A��0NSs���ID�I�WRK�^�� V��WV_]���> ��DI��q�@�{ /.�L_SE2�T���/�Z`��0��#�E_��u�v�j��SWJ�j� �Ȃ�	���=c�OH��z�PPJ�v�IR!��B� ��w�d��B8"����BASh���@ X ���V����?C�x�Q��RQDW��3MS���AX}�8�u�LIFE� �7�A1C�NJ���S��HӢ��Cs�>��C�`QN"�U��O�V� _�HE����S�UP�hbC�� _�Ԥ���_����[Q��Z��W���ו�Tb��XZ$ `1��Y2F�CM@T��t@��N�p�2r��9A �`�P.�HE��SCIZy֥�u��BN�poUFFI���p � �Q/40�<2671��wMSW9B 8�KEYIMAG�CTM@A��A�Jr|�0�OCVIET�N��C ��V L�t<���s?� 	�!� j:D�"pST�!x�0�� 0��Ѡ���0���EMAIL����@���ba_FA�UL��EH�CC�OU�p}$T@��F�< $���eS�]���ITvBUF@��q���T  ���	BdC�t����#��SAVb$)�e� �A� }���Pi�e@U�b`_ H���	#OT{BH�lcPր(0�
{��AX1#��X @��_GJ�
pP�YN_�� Gj�D��U/0e��M��*��T8�F��ِ�A!H�(@u��&�C_r@�@K�D����=pR���ugDSP �uPC�IMb��J����U��ЁEƀ��IP��su��D  �T!H0�c��TuA��HSDI�ABSC�ts��0Vzp*} ��$�#��NVW�G �#�$0� FJ�/ad�j�ASC��U�MER��uF�BCMP��tET�H�!AI��FU��D�U �a�@;⠂CD��O � ���R_N�OAUTg` J���Pp2��n4ĥPUSm5CF }5CI��.��k3� =K/H *}1Lp�� �Q��&�I���4#Q �6s��6ѡ�60��6��*�67�98�99�:J�T�8�:1J1J1JU1+J18J1EJ1RJ�1_J2mJ2�;J2�J2J2+J28J2�EJ2RJ2_J3mJ3�:3KJ3J/�G�8J3EJ3RJ3_J4�mB2qEXT�>aLC`��F�fF�5Q�9g�5 �FD�R�MT��V�C��C�wa}"C�RE�M,�FAj�OVM���eA�iTROVf�iDTm �jMX�l�IN�i���j�IN�D�`!�
xp /$DG���`opS�r9�D��`RIV)0�Qbj�GEAR�I%O0�K�bu�Nj�x��.؎��p�qj�Z_�MCM>�C�d`��U�R)2N ,{1��?g ��
 ?�p.I�?�qE���q��1T0lbO����P� �RIT5���UP2_ P Ѡ#TD= ��C�����qP�J�F .�BAC;Q T��$9 O�-)��OG��%E��3e&0IFI��e0X�0����PT���MR2ieR ivbY�vbLIq ��{g����f���J�b_mAN~F�_F��I4+�M;v`r}DG�CLF��DGDY&��LD�q>t5[�5�S�كk�S��M�� T�FS� l�T� P�)���
�/�$EX_)�@�)�1P�� ��*�3b�5b�s�G�!ieU � p�&2SWKO��DE�BUG�S��0�GRtY�zU�#BKU� �O1�@ O�P�O8��Π0��ΠM�S]�OO��SM�]�Eq�1pQ`_E� V $�X�� �TERM2�W�;�YTE�ORI�Ā6�X;���SM_ȗ�$7�Y;�ܰ�T�Ay�Zk�UPB�[�� -��QbV�$G���W$SEG�źאELTO���$USE0NFI����p����`���X$UFR����q00豈�D5h�OT1Ǵ �TA_ �C�NST�d�PATT!��Y�P'THJ!B0En�K0�ART� ����8����REL��&SHFTF"�_���_SH��M�!B0x�� ��n���Z���OsVR
#&SHI��ꅔU�2 �AYLO$ 5I1�_�8d���d�ERV�0*� } ��b?�d��Q�����A��RC
���A�SYMh���WJ�apE�����f�2�U��d�5����D5£�P#Gи!	�OR2d�M�h0GR!���\��΢�^�����k�] �E�.��TOC�졳q��OP��N z�3&1ʜ��aO�a> RE��R�#&O0��`�e��R]���������e$PWRSpI�M��[�R_���VcISy�r���UD��t�� ^>�$�H����_ADDR
9fH$�Ga�z�s��i1R� =_ H8�S� ��S��C��C��CSE�a����HSO0��` $���_D`�v��PR��1wHTT� UTH��a ({0OBJE�1u���$9fLE�P�-=b � �*g!AB_qT���Sk�#DBG�LV5#KRL"�H�IT�BG0LO:���TEM4$�0�b������SS�p�4�JQUERY_FLA��f WYA���ec��� PU�"B�IO0��4G���H��HB �IO�LN~�d/0i�C^��$SL�� oPUT_�$���Pwp�rSLA�� e/2�����ӡ��r�IO F�_AS�f��$L��U���#�04�#0����,�HYOgN!v'$FI!UOP�g ` l!9f�b>$�`E&�!��P����'�!E&�"�&؁IP_�MEMBk0T 7h X IPz�v��"_#0v����0��pOc6�1w�DSP��' $FOCUSB�Gv���Jhfi �q 60S��JOG�nW2DIS�J7��O��$J8�97†I6!�2�77_L�ABQ����0�8�1A7PHI�pQ�3�7D+�J7JRA4`P��_KEYp {�KILMON�=j&`$XR =~0cWATCH_ ��DӘ�U1EL� �y�`B�k GpG�V8P�-ffBCTR��fB�5��LG|�l ���+h�"��LG_SIZ{Y��E
��F
 �FFD�HI�H�H� �F�HM��F�@���C5V 
�5V
 5V�@5VM�5W��`S)@S����@Nv1��mx � ��R��4a�PÀU�Qk�L�S�RDAU�UE�A I���R�PGH���� BOO~�n�� C-"2�ITpGcd��)&REC-j�SCRN)&DI2`#S��RG�����cl�!#��b�!S�a"Wkd!�T!#J{GM�gMNCH�"FN�2�fK�gPRG�iUF�h	��h�FWD�hHL/ySTP�jV�hĀ�h`�hRSgyH!�{&C�Es��!#���g�yUt�g�¬f|@6#2�bG�i4�PO�Jz�ZeEsM�w82�iEX.'TUI�eIP�cw��c���c���`�a�����s��Jg��KaNO{�ANA"貇�gVAI�0zCL��~��DCS_HI���������O����S�I)��S'��hIGAN�@��C�aT��n��DEV�wLL��L�Q6@BU𠔠oa@��T��$�GE�M'9nDdѢ��p�a@ЅC�!��O+S1��2��3��s�83�����q �T0v�-�絡.e�IDX����-fL�b�STm R�PY0����� p$E��C ���  ����� ��r L*</��Q(6����6�EN 6�Օ~Kc_ s Y���P$ dKaD� �M�C�Rt �T0C�LDPm ��TRQ�LI`��e0x�f�FAL>1��_����DUA���LD������ORGe0�r���WX������Y���V�O�u �� 	���uu���Si�Tx��00�ްS�}[�RCLMCi�����{�m[�C0MI���O�v d�Q6�R�Q�00�DSTB���Y� ��{a��A�X��@�� �EXC#ES��ԑ��M��w���¹�+���5x(��_A�ʊ �l����V�K|�y q\*�2��$MB�LIE��REQU�IR����O��D�EBU��L�M{�zW�.!��B��i�E��N,03Ѩ�{�R��RkHV�DCE��TIqN3 `!�TRSMw0�p�S�N�����s<�P�ST�  |h�L�OC9�RI� 9�E�X��A��:�����O�DAQo%}��$@�Q΂MF�A��_���p�C��P��S�UP���FX��I{GG�"~ �0� �MQ���v�5@� %����m ��m ���О6#DATA����E�� 1�NP" N��[ t�MDIFA)?�!��H����1!� �Q"ANSAW�a!ܑS�!D��)��H3Q�$� ?�CU�@V_ >0��&�LO�P$�=ұ���L2�����3V�RR2I5�O  ��QAX�� d$CALI���NUG�2gRsINp<$R�SW0��K�AB�C�D_J2SE�����_J3v
�p1SP�@6 ��P�p�3��\���B�J���P�O���IM��[�CSKP ��$�P�$J�Q[Q,6%%6%,'��_cAZW��h!EL��<���OCMP�����1X0RT�Q�#�11�c@�Y�1��(�0:�*Z�$SMG�p�����ERJ��C0IN� ACߒ�@�5�b��1�_B��542d���14X҆f>9DI~!��DH �t30���$Vlo�Y�$�a$�  ��A�<�.A�����H �$BE�Ly lH�ACCE�L?��8���0IR�C_R���AT<w�c�$PS �k�L͠yP D��0Gx�Q�FPATH�9�WG�3WG3&B��#�_@�2�@�AV���C;@��0_MG|a$D�D�A@[b$FW�(����3�E�3�2�HD}E�KPPABN.GROTSPEE�B���_x�,!��DEF�g��1͠$USE)_��Pz�C ����YP�0V� �YN���A{`uV�8uQM�OU�ANG�2�@O9LGC�TINC~����B�D���W���ENCS����A�2��@INk�I&Be���Z�, VE�P'b2�3_UI!<�9cLOWL3��pc x��UYfD�p��Y�� ��Ury�C$0 fMOS`�Ɛ�MO����V�PE�RCH  vcOV�$ �g9��c��\bYĀ���'�"_Ue@0��A&BuL������!epc�\jWvrfTRK�%h�AY�shчq&B��u�s���&l��Rx�MOM|���h�ﰞ �Ą�C�sYC���0D�U��BS_BCKLSH_C&B��P �f�`}S�7��RB��Q.%CLAL��b?�8�pX�t�CHKx�H��S�PRTY�����e�����_~��d_�UMl�ĉCу�ASsCLބ PLMT��_L�#��H�E ������E�H�`-��Q#p_��hPC�aB�hH��ЯEǅCw���XT�0�GCN_b(N�þ���SF�1�iV_RG�e�!��&B����CATΎSH ~�(�D�V��f�0'A�	� �@PA΄�R_Pͅ�s_y�뀎v`�`x��s����JG5��6Ф�G`OG���rTORQUQP��c�y��@�Ңb�q�@�_W �u�t�!�14��33��3�3�I;�II�I�3F��&������@VC"�00���©�1��2�8ÿ�¶�JRK�����綒 DBL_SMt�QO�Mm�_DL�1O�GRV:�3ĝ33��3�H_��Z@a��COSn˛ n�LN ���˲��ĝ0��� �� e��ʽ̃��Z���f��MY���z�TH|��.�THET0beNK23�3Xҗ3��[CB]�CB�3C��AS���e��ѝ3���]�SB�3��h�GT	S@! QC���'y�x�'����$DU�� ;w	��Q�����q9Q����$NE$T�!I�����)I7${0LсAP�y��`�k�k�LCPHn�W�1eW�S�� �������W���������{0V��V��0��UV��V��V��V��UV��V�V�H��@����7�����H��UH��H��H�H��O��O��OF	��O���O��O��O��O*��O�O��FW�}���	�����SPBA�LANCE�{�LmE��H_P�SP1��1��1��PFULC5\D\��:{1��!UTO_���ĥT1T2��22N���2, ����q^P<�-B#�qTHpO~ |�1$�INSEG�2�{aREV�{`aD3IFquC91�('o21�dpOB!d�=���w2��7P���LC�HWARR�2AB����u$MECH`��ДQ�!��AX�q�PB��&r�~2�� �
�"��1eROBF�`CR r�%��S0�MSK_�4� WP �_OPR�1�2(47Qst1�,`*R`(0)cB�(0|!IN!��MTCOM_�C���0�  ��@0 �A$NOR�Ec�2�l ~2�� 4�GR��%F�LA!$XYZ�_DA��LP;@DE�BU�2 �0lR�0�u ($mQCODS�G �2�r� �p�$BUFIND�X*P0;@MOR3� H%0�p�0���:@�p�QB�"�1c��NF�TA9Q�"@�2�rG.B� �� $SIMUL����0�As�AsOB�JE3�FADJUyS�H�@AY_I��:xD�GOUTΠ�4��p�P_FI�Q=8AT#�Y,`W�1P @+�PQ+ 9�uDjP�FRI �PUT0�R�O�
`E+�Sp�O�PWO��0�,>@SYSBUi� @$SOP�QBy��ZyU�[+ PRUNn2�UPA;0D�V�"�Q��`_�@F��PP!ABx�!H��@IMAGS�i%0?�P!IMQA�dIN$��RcRGOVRDEQ�R�@�QaP�Pc�� L_�0�feÂސRBߐ<p}X�MC_ED'@*�  H�Ni M�bG��MY19F�0Ea�SL30� x �$OVSL�S;DIsPDEXǓ�fH֓Hq�bV+��eN�a 
��Pp�cwx�bw�=�d_SET�0�� @�Cr�%9�R)I�A3�
Vv_��bw�{qnq0-!�@� ��4BT� àAT�US�$TRCpA�@PB�sBTM�w�qI�Q�d4F��s�`.0� D%0E�P�b�rr�E1"�qQpd��qEXE�p���a��"��tKs�Rp&0�pU�P�01�$Q `X�NN�w���d���y ��PG|5� $SUB�q�%xq��q|sJMPWAI2$�Ps��LO ��1�
 �E$RCVFAIL_C@1�PÁR%P�0�#���Ȕ� ��
�R_PL|sD�BTBá���PBW�D��0UM��I�G�Q `�,�TNL ��b�ReQ�2���qP��@EǓ��֒���DEFSP� �� L%0� ��_8���CƓUNI�S�w�Đe�R)��+�_L�
 P�q�qPH_�PK�5��2RETRIE|s�2�R{B����FI�2� � �$�@� 2���0DBGLV�LOGSIZ�C� ����U�"|�D?�g�_)T:��!M�@C
 #�EM��R��y0�8C�HECKS�B�Po01��0.�0R!:LbNMKET��@��3�PV�1� -h�`ARp� �1)P��2>�S�@OR|sF�ORMAT�L�C!O�`q����$Z���UX�P!r�LI|G�1�  ˣ�SWIm �a1A�X,�G�AL_ G� $`@��B�a��CS2D�Q$E�1��J3DƸ�{ T�`PDCK�`|�!LbCO_J3�����T1׿� ��˰C_Q�` �; ��PAY��S2�u�_1|�2|�ȰJ�3�ИˈŬƗ�tQTWIA4��5��6S2MOMK@��������4��y0B׀AD���������PU��NR ��C���C������4��` I$PI N�u�41�žӁ�:q� R~ȇ��ٯ��:�h� �a�֬��ց�1�'|1R\uSPEED G��0�؅��7浔؅ �%P7�m�F��U��؅SAM =G��7眪�؅MOV	B�  e0�� ��c2��v��� ���� ���c2nPsR�����İ$QH���IN 8�İ��?�[�6�؂A����X����GAMM��q�4$GETH1R@�SDe�mB
�OLIBR[�y�I�7$HI�0_5a@c2E`@#A@ 1LW^U@	�1a¬&o�ʱC=�n S`ރp �I_ ��pPmDòv�ñ'�����mD��	ȳ {�$�� 1��0IzpR� DT#|"c���~ LE^141�qw�a�?�|�MSWFuL�MȰSCRk�7�0��Ѻv���Z 0�P�@9@����2�cS_SAVEc_Dkd%]�NOe�C�q^�f� ��uϟ� }ɕQ��}���}*m+��9��ժ(��D�@���� �������b31�RA�Mam�7
5�#��^�����Mtա � �YL��
A'�VAS	BtRna`7GP �B
Bl3
A%`�GSB1W? �2�2cЬ3doBB1M&@�;CL�8����G�b�1v���M!Lr� �N�X0�d$W @�ej@b��  @=�BD�BK�B� -�> �P����ycİ%X �OL�ñZ�E����uԣ ��OM�R/d/v/�/�/P��A�j	�Le�_��� |��H ��jV ��yV��yP�ʗW�V�ʡE���FZ��8�t��NTP=��PMp�QU�� � 8�TpQCOU,�Q�THQ�HOY2`H�YSa�ES��aU�E `"#�O��� �  �P�0�rUN��p�3��O$�J0� P�p^e������OOGRA�qk22�O�d^eITm�aB`/INFOI1���k��ak2��OI�b�{ (!SLEQ(� �a��`�foaS� ���� 4TpENA�BLBbpPTION�|s����Yw��1sGCuF��O�$J�,ñfb���R�x!��]ot�ROS_ED�ŀJ0� �N��@K��᪃ES NU��w�xAUT,!�uCOPY�����v�8 �MN���PR�UT�� �N�pOU��$Gcbn��R_RGADJI1�2�3X_B0ݒ$ ����@��W��P������@㊀��EX�YCZLB��NS6u�N0άLGO�A�NY�Q_FREQZ�W`���+�p�\cLAm�"����Ì�uCRE�  c� IF�ѝcNmA��%i�_GmSTATUQPmMAIL�� 1��y�d����!��ELE�M�� �7 DxFEASIGq2��v���q!�er$�  I �`�"��ae�|I��ABUq�E�`D�V֑a�BAS��b� �[�Ub�r % $�y���RMS_TR C�ñj���Ca��ϑ���,r���C�YP	~ � 2� g� �DU�����Ԣ�0-��1��1���qDOUd�ceNrs��PR30z;p�rGRID�a�UsBARS(�TY�Hs��OTO�I1��P`_��!ƀ��l��O�@7t� � �`�@POR�cճ��.ֲSRV��)���DI. T���!���+��+�4)�5)�6J)�7)�8��aF���:q�M`$VALAU|�%� 0>1F6u�� Cu'!�ab���� (gpAN#ĳ�R�p0� 1TO�TAL��[��PW��It�&�REGEN$�9��SX��sc0��Q���PTR��Z�$�C_S ��9дsV���t���rb�E��x�ap�"^b�p��V_H���DA�C����S_Yh4!�B<�S�AR�@�2� f�IG_CSEc���˕_b`F��C_����w��?rp��%�b�H�SLG#�
I1��p"=���4d��S�2̔DE�aU!Tf.p��TE�@>���� !a����Jv�,"��IL_�MK��z�н@TQ@�P�a����2VF�ECT�P���^�Mu�[V1t�V1��2��U2��3��3��4��4����С���1�"IN	VIB�@N�; �!B2>2�J3>3J4>4�JI05���"���=p�MC_F`3 � L!!�r��M= I��M� �[PR�� KEEP_HNADD��!f�C�A�� !����"O�Q �I����"��?�"REM9!�ϲ^�uzU��e!HP�WD  S/BMSKG�a	!�B2B�
#COLLAB�!��2����4�o��`IT��A`��D� ,pF�LI@��$SYNT� ;,M�@C>��%пUP_DLYI1�MbDELAm ј��Y�PAD�A<2QSwKIPE5� ��``On@NT�1� P_``�b�'�`�B]0 �'���)3��)��)O� �*\��*i��*v��*��z�*9�J2R�*���?sX��T%�|1�{2ܐ�|1�a���`RDC!F� ���pR�sR�PM�'R�^��:b�2�RGEp�p2��3d�FLG�Q8�J�t�SPC�c��UM_|0��2TH�2NP�F@o0 o1� �0EF�p;11��� l[P�E-Ds#ATWo�[� w�B�`�d�A�p3�B�fcAHnP�B��_D2gB�mOO�O�O�O�O
�G3gB��O�O_ _(2_D_�G4gB�g_y_��_�_�_�_�G5gBĀ�_�_oo,o>o�G6gB�aoso�o�o�o�oW _D7gB��o@�o&8�G8gB�[m����E)S����\@ǡ`C�N�@�_@wE���^� @o��m�I�O�ፉI�ޡj�P�OWE!� �W�: �1���0� y�5%Ȃ$DSB;����֒ �h CL@��ެ1S232s�� Ɍ�0�u.��IC3EU{���PEV@�џPARIT�њ�O�PB ��FLOW�TR2�҆]����CUN�M�UXT�A���INTER�FAC3�fU���i�SCH�� �t� � ˠE�A$L����OM��A�0"נI���/�A�	TN���Tо ��ߓ��EFA� �"!�Ҏ��� u!��� �O�� &*�� ������  2� ��S�0�`�	�' �$3@}%:B��䎣�_���DSP���JOG��V�h�_P�!s�ONq0%�0����K��_MIR����w�MT7��A�P)�w�>@"���;AS�������;APG7�BRKH����G �µ!! ^���i���P���<����BSOC��w�N���16�SV�GDE_OP%�FSPD_OVR��u �DвӣOR$޷�pN��߶F_���6��OV��SF�<���
�F0����UF�RAF�TOd�LC1Hk"%�OVϴ ��W[ ���8�Ң��͠;�  @ BT�IN����$OFeS��CK��WD����������r���TRr��T�_FD�� �MB_C �B��B����(�.Ѻ�SVe��琄�}#��G)�<�AM��B_0��jթ�_M@�~�x�ቂ��T$CA�����De���HBKX�����IO�������PPA���������Տթ���DVC_DB��?����A���,�X� b��X�3�`���3Z0����ϱU8󳠈�CAB�0��ˠ��c� �Ow�U�X��SUBCPU�ˠS�0�0�R�����!�A�R�ł�!$HW_Cg@A��!���F��!�p� � �$�U r�l�e�AT�TRI��y�ˠCY�C����CA���FLT ��������vALP׫CHK�o_SCT��F_e�cF_o����FS�J�j�CHA�1��98I�s�8RSD_!�0���恩�_Tg�7��� �i�EM,��0M"f�T&� @�&�#ޮDIAG��RAOILACN���M�0 �"��1���L���{�PRB�S   ���C4�&�	��F�UNC�"��RI	N�0 "$�7h�� S_��(@��`�0p��`A��CBL� �u�A����D�Ap�a���LD@ܐð�����j���TI%��@�$CE_RIAAV��AF�P=�>#,��D%T2� C��a��;�OIp��DF_aLc�X��@�LML��FA��HRDYO,���RG�HZ 7�����%MULSE�� �����k$J�ۺJ����FAN?_ALMLV�1�WRN5HARD�r��Fk2$SHADOW|�Gq��O2 s�0N�r�J�_}����AU- R+�TO_SBR���3���:�e�6�?�3MPIN�F@{��4��3R3EG�N1DG�6C1V��s
�FLW��}m�DAL_NӀ:����B�	����a�vU�$�$Y_B�ґ u�_�z��7� �/�EGe����ð�AAR������2p�G�<�AXE��wROB��RED���WR��c�_�M��S�Y`��Ae�VSWWcRI���FE�STՀP����d��Eg�)�$�D-�{2��BUP��t\V��D��OTO�19)���ARY���R0���<rנFIE����$LINK�!GkTH�R�T_RS���E��QXYZt��Z5�VOFF��b�R�R�X�OB���,8d����9cF�I��Rg��􃻴,��_J$�F�貿S��q0kTu[6��1�w �ad�"�bCԀ+�DU�º�F7�TUR0X#�e�Q�2X$P�ЩgFL�Pd���@p�U�XZ8���� 1�J)�KʠM��F9�p��ӓORQ����fZW30�B�O Pd�,��t����A�t'OVE�q_BM���q ^C�udC�ujB�v�w0L�wg��tAN=�Q �qD!`A�q��=�}��q �u�q���dC��"���SERϡj	�E��HT�ńAs�@�Ue�X��W����AX ��F����N�R�� +��!+�� *�`*��`�*��`*�Rp*�xp*�1 �p*�� '�� 7�� G� � W�� g�� w�� ���� ��� ��đ��DEBU=�$8D3�h����RAB�����r�sV��<� 
�� i�`A��-񷧴���� ��a���a���a��Rq���xqJ$�`D"�R9cL�ABOb�u9�F�G�RO��b=<��B_���AT�I`�0`�����u���1��AND fp�ຄ���U���1ٷ ���0�Q�������PNT$0M�SE�RVE�y@� $�%`dAu�!9�PO��[0ЍP@�o@*��c�x@�  ]$]�TRQ�2
\�d�Bf��j�D"2�{��" � _ � l8"T�c6ERRub��I��VO`Z���TO	QY�V�L�@)�1R��J� G;�%�Q�2 [�T0e�� ,7�ř���]�RA#� 2'� d@����r�7 �Y@$�p��t ��OC�f���  ��COU�NTUQ�FZN_wCFGe�� 4B�F��Tf4;�~�\� ��
�ӭ�uC� ���M: �"`A��U��q: �FA1 d�?&�X�@=����_B�A<�����AP��o@HE�L@��� }5�`B_BAS�3�RSRF �CSHg�!��1
ש�2��U3��4��5��6���7��8
ל�ROO0�йP�PNLdA�c�ABH�� ��ACK���INn�T��GB$�Uq0� +\�_PUX��@0��OUJ�PH�H���, u��TPFWD_KAR��L@��REGĨ P�P��]QUEJRO �p�`2r>0o1I0������P����6�QSE�M��O��� A�S�TYk�SO: �4D�Iw�E���r!_�TM7CMANRQܨ�PEND�t$�KEYSWITCaH���� HE�`�BEATMW3PE��@LE��]|� U���F>��S�DO/_HOMB O>�_�EF��PR>a9B�ABPx�CO�!��#яOV_M�b[0# I�OCM�d'eQ�ъ�HKxA� DH�QG��Ue2M�x����cFORCC�WAR�"�Ҋ�OM>�@ � @r�:#��0UHSP�@1&2*&&3&&4�A��sЕO��L"�,�HU�NLO��c4j$E�Dt1  �SN�PX_AS��� �0+@ @��W1$S{IZ�1$VA��~�MULTIPL���#! A!� � $��� NS`��BS�ӂAC���&F'RIF�n�S��)�R� NF�ODB�U$P���%B3=9G��Ѫ�y@� x��S�I��TE3s�r�cSKGL�1T�R$p&���3a�P�0STMTd1q�3P�@5VBW�p��4SHOW�5���SV��_G��� Rp$PCi�oз��kFB�PHSP' 1Av�Eo@VD�0vC��� ���A00޴RB% ZG/ ZG9 �ZGC ZG5XI6XI7�XI8XI9XIAXIB�XI ZG3�[F8PZGFPXH��XdI1qI1~IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1 Y1Y1YU2WI2dI2qI2~I2�I2�I�`�X�IQpT�X�I2�I2�I2�I2 Y2Y2Y�p�h�dI3qI3~I3�I3��I3�I3�I3�I3��I3�I3�I3�I3� Y3Y3Y4WI4�dI4qI4~I4�I4��I4�I4�I4�I4��I4�I4�I4�I4� Y4Y4Y5�y5�dI5qI5~I5�I5��I5�I5�I5�I5��I5�I5�I5�I5� Y5Y5Y6�y6�dI6qI6~I6�I6��I6�I6�I6�I6��I6�I6�I6�I6� Y6Y6Y7�y7�dI7qI7~I7�I7��I7�I7�I7�I7��I7�I7�I7�I7j Y7Y7T >A�P� Uc�� �l�נ��
>A820��j���RCM2����MT�R��|���Q_��R-��ń�����[�YSL�1�� � �%^2��-4�'�4��-Y�BVALAU�Ձ���)���FJ��ID_L���HIr��I��LE_������$OE�SA~b�� h 7�VE_BLCK�¡1'�D_CPU 7ɩ 7ɝ �����E����R � � PW��>�%0��LA�1Saѝî����RUN_FLG �Ŝ������ �����Ą����H���Чī�TBC2��_� � _ B���� br� W?�eTDC����X��3f�S�THe������R>�k�ESERV!EX��e��3�2 ��d��� �X ;-$��LENX�Ԙe�Ѕ�RA��3�L'OW_7�d�1��ҴM2 �MO/�s%S80t�I��"�ޱH�����]�DEm�41LACE�2�CCr#"�_MA� l��|��GTCV����|�T� ������0Bk�)A�|�)AJ��%EM7���JH��B@k�X�|��с2p �0:@q�j�x JK��VKX������ы�J0����JJv��JJ��AAL��P�������4��5��� N1�� ����%LF�_�1� Ҡ лCF�"� `�G�ROU���1�AN�6�C�#\ REQUsIR��4EBU�#���8�$Tm�2�����|ё %�� �\�APPR� C�A�
$OPEN��CLOS<�S�v��	k�
��&� �<�MhЫ���v"/'_MG�9CD@�pC ��DBRKB�NOLDB�0RT�MO_7ӈr3J��P������ ��������6��1�@ p0�%��� � ����'��-#PATH )'B!8#B!�>#� � 9�@�1SCA��l�8IN��UCL�]1� C2@UM�(Y "��#�"�����*���*���� PAYLOA�J2LڠR_A	N`�3L��9
1�)�1CR_F2LSHi2D4LO4�!H7��#V7�#ACRL_@�%�0�'�$��H����$HC�2FL�EX�;J#�� P�4�F߭߿��|�0��� :�� ��|�HG_D����|���'�F1_A�E�G6�@H�Z�l�~���BE�� �����������*� �X�T,�C���@�XK��]�o�^Av�T&g�QX >�?��4TX���eoX �������������������	-	"J@� �/�M_q~�۠cAT�F�6�ELHP�Ѭs�J� � J�EoCTR�!�AT�N���v|HAND_VB��1��$7� $:`F2Cx�-��SW�A"�� $$M,0 0�_Y�ni��P\����A��� 3�����<AM��_AmA�|��NP�_DmD�|P\ G��E�ST�aM�nM�NDY ��� C����0��>7 _A>7Y1�'��d�@i`�P��������":J$�� �O�4D'"r�J���A'SYMl%A�� l&!��@�-Y1�/_�}8 � �$��� ��/�/�/�/3J	<�:;�1�\:9�D_VI�x�|��V_UNI�����cF1J����䕶� Y<��p5Ǵ�y=6��9 ��?�?>�wc�4�3ߩ�$� AS�S  ����s�  �{�h�VE�RSIONp��=��
��IR�TU<�qσ�AAV�M_WRK 2 ��� 0  �5z��������� ��	8�)�L�{����:�w�^�|�(ܛݧ��7ѭ���������BSwPOS� 1��� <�� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������//�1/C/U/ⰑAXL�MT��X#�%�  dj$INs/�!i$PRE_EXE�(A� �&)0�q��������LARMRECOV �ɥ"
�LMDG �����[/LM_IF �ˆ!X/c?u? �?�?�:Q?�?�?�? OM, 
0�8O�4��cOuO�O�O�NG?TOL  ��ЏA   �O�K��P�P)�O ;� ?6_,_>_P_{� $BR_�_w�o_�_�_ �_�_�_o�_'oo7o]o�!��O�o�o�o�o �o�o�o+=O�a�PPLICA�T��?��� ��J`Hand�lingTool� �u 
V8.?30P/33�@lt���
883�40�slu
�
F0�q�z{�
�2026�tlu���_�7gDC3�pJ  �s�Nonelx� �FRA�������B�TIV�%�s�#��UTO�MOD� E�)P�_CHGAPON������ҀOUPL�ED 1��� ���"�4�uz_CUREQ 1��S  � >�>�*����4��!��x��~� ��u���Hm����HTTHKY����w���7� ���%�C�I�[�m�� ������ǯٯ3���� !�?�E�W�i�{����� ��ÿտ/�����;� A�S�e�wωϛϭϿ� ��+�����7�=�O� a�s߅ߗߩ߻���'� ����3�9�K�]�o� �������#����� �/�5�G�Y�k�}��� ����������+ 1CUgy��� ���	'-? Qcu����/ ��/#/)/;/M/_/ q/�/�/�/�/?�/�/ ??%?7?I?[?m??���P�TO�@����DO_CLEAN܏|��CNM  �K >�aOsO�O�O��OD�DSPDRY�RO̅HI��=M@ NO_'_9_K_]_o_�_��_�_�_�_�_�_J�MAX�p�4�1���a�X�4"��"���PL�UGG���7���P�RC�@B;@?K�_�_ebOjb�O��SEGFӀK�o�g�a ;OMO'9K]�o�aLAP�O~Ǔ� ������/�A��S�e�w���΃TOT�AL-fVi΃USE+NU�`�� ������P�RGDISPWMMC�`{qC�a&a@@}r��O�@f��e��_STRI�NG 1	ˋ
��MĀS���
`�_ITEM1j�  n�������� ��Ο�����(�:� L�^�p���������ʯ�ܯI/O S�IGNALd��Tryout M�odek�Inp��Simulat{edo�Out.�OVERR�@� = 100n�In cycl"��o�Prog A�bor8�o��S�tatusm�	H�eartbeat�i�MH Fauyl����Aler�� �ݿ���%�7�I�8[�m�� �3f� �1x����������� *�<�N�`�r߄ߖߨ߀�����������WOR�`f�L���&�t� ������������ �(�:�L�^�p�����8������POd��� ��d���%7I[ m������ �!3EWi��DEV����� ���//'/9/K/ ]/o/�/�/�/�/�/�/��/�/?PALT ��81d�?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O&?GRI`f��AP?�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHo�OR�̀a �OZo�o�o�o�o�o &8J\n��������noPREG<>%��o�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~������$ARG_�L�D ?	����ӑ� � 	$�	+[�]�����ƐSBN_CON?FIG 
ӛ&��%� �CII_SAVE  ��E�<�ƐTCEL�LSETUP �Ӛ%  OME�_IO��%M�OV_H������R�EP�l���UTO�BACKt�0��FRA:\�c ���_�'`����=�� J� 	������ͿpĿֿ�6����	� 1�C�U�g�yϋ��� ����������ߜ�5� G�Y�k�}ߏߡ�,��� ���������C�U��g�y����a� � )�_�_\AT�BCKCTL.T�MP DATE.D;<��	��-�?���INI;0p�8�~�MESSAGT��^�_�ېi�ODE_AD��W�8�H���O�����PAUS��!��ӛ ((O ֒��
��*N< r`��������"����TSK�  ��=�C�	�UgPDT��\�d����XWZD_ENqB\�4��STA[��ӑ�őXIS&�U�NT 2ӕ`� � 	S
/�� 2//V/A/z/e/�/�/��/�/�MET�`2�P�/?�/<?�)�SCRDCFG }1C`�	�\�\�1?�?�?�? �?�?�?6��QX��? ?OQOcOuO�O�O O�O $O�O�O__)_;_�O�O���GR�����zS��NA��қ	��wV_EDZ�1�e9� 
 �%{-��EDT-h_0ʪ�_o�`/A���Q-��_�	���x���_�o  ���e2�oɫko�o�6k�o@!hozo�o�c3Y �o��o�n��4F�j�c4%��r�� �nN��� ����6��c5�a�>����n��� ̏ޏt���c6��-� 
�Q��n�Q�����@�Ο�c7����֯��n����d�v�����c80U��_����0
 }~�@�0�B�ؿf��c9!���nϵ� }Jϵ���0Ϥ�2φaCR�oį 9�K���������n����zP�PNO_DE�L�_xRGE_UN�USE�_vTIGALLOW 1�Y�~�(*SY�STEM* 3	�$SERV_GRp�R 69���REGB��$d� <9�NUMxg��z�PMU��> 5LAY�  <�PMPAL|[��CYC10�����������ULS�U��{�����D�L��N�BOXORI�k�CUR_;�z��PMCNV���;�10���T4DCLI�4�V���� ���'9K]�oR�zPLAL_OUT Dcc�QWD_ABOR���	��ITR_RT�N���Y� NON�S8� �CE�_RIA_I�j�<F_1���B =[_PARAMGP 1�w`_�����Cp  .�� � � � �� � � � Ҫ � � � �7  D5`D$3!�g-�<$�H$�T$�� DX � �X "� B�D1� 9�X @� 6?� <H=E��ONFIy��n�!G_P��1� �e�U??0?�B?T?f?x?�?�!KP7AUSX�1�UR ,Z��?�?�?�? �?OOOTO>OxObO �O�O�O�O�O�O_�2�O_ey�PCOLLECT__a�Y5auGWEN��pI�"cR QNDEOS��W��1�234567890�W�S�u�_�Vy'
 H�y)�_#o S��_ohoT�AoSo�o wo�o�o�o�o�o�o< +�Oas� �������\��'�9�K���o��VQ�2�W[ � t�VI�O �YcQy�H&�8�J�\��TR��2؍(��
��j��  ����%^�_MOR҂!�� + �'� 	  �5�#�Y�G�}�k���D�Ӂ"��2?�!��!3 ҡ�Kڤ�
�$R_#*_	���C4  AS yC � x�A3!z � BC!�PB/!�PCo  @*�����:d�
�I�PS$���T��FPROG %�*6߼�8��I����&�RҴKEY_TB�L  )VR�� �	
��� !"#$%&'�()*+,-./��W:;<=>?@�ABC��GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~��������������������������������������������������������������������������������͓���������������������������������耇���������������������9��1��LCKۼ3����STA�д_WAUT��O(���U�INDtTD�FQRg_T1_�Q�T2�߰7$����XC� �2����P8
S�ONY XC-5�6������@����u� ���w��HR5���cT0�B�7T�f�ACffrꬿ���� �� �����5�G�"�k�}� X��������������ǼTRL��LE�TEG��T_S�CREEN ~�*kcsc:�U$MMENU �1&�)  <���y�� Ã�=&sJ \������� '/�/]/4/F/l/�/ |/�/�/�/�/?�/�/  ?Y?0?B?�?f?x?�? �?�?�?O�?�?COO ,OyOPObO�O�O�O�O �O�O�O-___<_u_ L_^_�_�_�_�_�_�_ �_)o oo_o6oHo�o lo~o�o�o�o�o�o �oI 2X�hz����� _MANU3AL�ߕ�DB���L+�DBG_ER�RL��'��C �\�n�����NUMLIMK��d �p�DBPXWORK 1(�I�ޏ����&�Ž�DBTB_@ Q)�������qDB_AWAY��_�GCP  �=s�װ�~�_AL��D�z��Y��M � ��_)� 1*�
���
͏����l6�@�_M{�ISA��@B�P�ONTImMJ� ��p��ƙ
�ۓMOTN�END߿ڔREC�ORD 10}�� �>�?�G�O� ���?���2�D�V�h� ��p������*�߿� Ϛ���9Ϩ�]�̿�� �ϥϷ�R���J���n� #�5�G�Y���}��ϡ� ���������j��� C��g�y������ 0���T�	��-�?��� c���\���������� P�����;��_q �����(�L %�4[�� ���^t�l!/ �E/W/i/{//�// �/2/�/�/??�/z��TOLERENC懔B�В��L����CSS_CNS�TCY 116�  ?Β�?�?�? �?�?�?�?OO&O8O JO`OnO�O�O�O�O�O��Oc4DEVICEw 126� b� *_?_Q_c_u_�_�_�_�_�_�_?�d3HND�GD 36�C}z�^LS 24]�__oqo�o�o�o�o��o�_e2PARAM� 5�B��t�d�c4SLAVE �66�e_CFG �7��gdM�C:\e0L%04�d.CSV�o��c�|�r�"A �sCH�p&a&��n��w��f�r�����ÀJP�>��\_�CRC_OUT �8U����oEpSGN 9U�Ƣ�02-OCT�-22 14:4�1�p����9V UBu1�݁�nހ���\�o��I�m��P�uG���@uVERSIO�N ��V�3.5.11E�E�FLOGIC 1�:ݫ 	6���|�C���^�PROG_ENB����͢.��ULS{� ���^�_ACCLIM^|��Xs��?WRSTJN[���ţ�^�MO��¡Zr�,�INIT ;�ݪs5� *�OP�T$p ?	i�B�
� 	R575��c��74��6��7F��50��R�Ƣ2���6��X�y�TO  ����?�Y�VP�DKEX�d#��@W�PATH A���A\E�����7;I�AG_GRP 2�@�k,�"	 �E�  F?h� Fx E?`�D��û��V1"��ü��T0K�9�Cf��py�pY�dC��pq�B�i��ùmp4m5� 7890123�456��;���� � A�ffA��=qAةpхA��HAĩp��������Ac��Mk���@��t�p�p��W0A�T0T0�pB4ü Qô����
���(�A���A�
=A��L���A��
�A�Q�A��������e������e� Pe�:��{A��d�����dѩp�������A���������r߄ߖߨ�|��@�EG�A@�p_:�RA5d�/��U)��#P�d�l�������"�4�F�@�POz�AJ��c�?���9p�A3\)A_,��A&�����0��������@�c�P�]��AW�P��J��C��<d�4:�-d�%G��(� :�L�^�@���$ HZ��.|��� �bt� 2V h�xm�����[����s�����=�
=�=�G��>������7���8���b�7�7��%�@ʏ\"&��p�.%��@�Ah�p9 A��<i���<xn;=R��=s��=x<��=�~Z�;���%<'�'�~� �?+ƨC��  <(�U�� 4"����&�C���%ùf��@?� �?�?@?R?g��$ ^?�?"?�?�?�?�?�?��?)7L?S��FB$�/"Eͽ,�>OG�ΐԬq���sD�L4�x�CA��Gb�tφ���-_7_�C��_;�/_�N�ED  E�  �Eh� D[PbRpD_¿�_�86� �_�_
z{_�_w_o�K:o@bùQm)o�o�o�o�o�o�o�o ɼC�T_CONFIG; ��Yt؃�eg��ԱSTBF_TTS��
ęVs3���
�iv�[�MAU���Y�M_SW_CF*pB��  �Q�OCVI�EW}pC�}����_�!�3�E�W�i� ;��������ȏڏ� {��"�4�F�X�j��� ������ğ֟����� �0�B�T�f�x���� ����ү������,� >�P�b�t�������� ο��ϓ�(�:�Lϰ^�pς��|RC�sDJ�r!ϐκ��������7�&�[�otSB�L_FAULT �E���xu�GPM�SK_w��pTDI�AG F.y�q��IUD1: �67890123#45��;x�MP�o!� 3�E�W�i�{���� ����������/�A�F�X W!�J�"
�|��vTRECP����
�����M� (:L^p��� ���� $6�]�o�l��UMP_?OPTION_p��F�TR�r`s����PME^u�Y_T�EMP  Èϓ3B�pp �A  �UNI�pau!��vYN_BRK �G�y��EMGDI_STA%�1!�G%NCS#1H�{ ��K��9�/_}d d�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO� �O�O�O�O�I�!�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXo�JO�o�o �o�o�O�o�o+ =Oas���� �����'�9�K� ]�wo���������oۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�o�]��� ����ɏ�����	�� -�?�Q�c�u������� ��Ͽ����)�;� M�g�y��ϕϧ�]�ӯ ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�_�q�{� ������������� �/�A�S�e�w����� ����������+ =Oi�s����� ���'9K ]o������ ��/#/5/G/ak/ }/�/�/��/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OY/KOuO�O�O�/ �/�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oQOcO moo�o�o�O�o�o�o �o!3EWi{ �������� �/��o[oe�w����� �o��я�����+� =�O�a�s��������� ͟ߟ���'�9�S� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�K�9�g�yϋ� ������������	�� -�?�Q�c�u߇ߙ߫� ����������)�C� U�_�q��9�Ϲ��� ������%�7�I�[� m�������������� ��!;�M�Wi{ ������� /ASew�� �����//+/ EO/a/s/�/��/�/ �/�/�/??'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O=/GOYOkO }O�/�O�O�O�O�O�O __1_C_U_g_y_�_ �_�_�_�_�_�_	oo 5O'oQocouo�O�O�o �o�o�o�o); M_q����� ����-o?oI�[� m���o����Ǐُ� ���!�3�E�W�i�{� ������ß՟���� ��7�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���/�9�K� ]�oω��ϥϷ����� �����#�5�G�Y�k� }ߏߡ߳��������� �'��C�U�g��w� �����������	�� -�?�Q�c�u������� ���������1�; M_����� ��%7I[ m������ �)3/E/W/i/� �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?O!/+O =OOOaO{/�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_O#o5oGoYosO eo�o�o�o�o�o�o�o 1CUgy� ������o� -�?�Q�ko}o������ ��Ϗ����)�;� M�_�q���������˟ ݟ�	��%�7�I�[� u��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ�a�� �/�A�S�m�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� e�o��������� �����#�5�G�Y�k� }�������������� ��1C]�Sy� ������	 -?Qcu�������� �$E�NETMODE �1I^��    �(/:+
 RROR�_PROG %�*%}/�)X%TA�BLE  +�h�/�/�/�'X"SE�V_NUM &"?  �!!0�X!_AUTO_ENB  D%#U$w_NO21 J+�9!2  *�*u0�u0�u0�u0(0�+t0�?�?�?N4HI�S3
 G;_AL�M 1K+ �2u< +�?/O@AOSOeOwO�O�?_2.T0  +s1:"��J
 TCP_VE/R !*!u/�O�$EXTLOG_7REQ�6�E9 S�SIZ)_TSTK�FYc5�RTOoL  
Dz�2��A T_BW�D�@�P<6�Q8W_D�I�Q L^�G48$
?"�VSTE�P�_�_
 �POP_�DOh_!FDR_?GRP 1M)B1�d 	�Ofo: W`��������glpw��qŗ��I ����fWc�o�m�o �o�o�o(L7�I�m��zA�f��A�ز>����� 
 E��	�q�@(�C���<�'�`�K�C`}d�C��N��B�y{��F�@UUT��UTF�Ϗj��s���s�OHcEP]���O��#M���*�KA����?��pF��:6:�N�r�9-��z�������������+FEAT?URE N^�P�>!Han�dlingToo�l � mpBo�Englis�h Dictio�nary�
P�R4D St�ڐard�  o�x, Analog I/O��  ct\b+�g�le Shift��  !*�uto� Softwar�e Update�  fd -c�m�atic Bac�kup�IF O���groun?d Editސ��g R6Ca�mera3�F7�P�art��nrRn�dIm���psh�i��ommon calib U����n����Moni�tor�CalM��tr�Reli�abL��RINT�Data Acquis�Z�Ϡ~C�iagnos���0�<�almC�oc�ument Vi�ewe�\���C�u�al Check Safety���  - B�Enh�anced Us抰Fr���8 R�5�xt. DI�O �fin� (��@ϲend��Er�r�Lm� D ph^���s	�EN��r.�հ �P�rd�sFCTN /Menu��v8����m�FTP InN'�facN�=�G���p Mask E�xc��gǱisp���HT^�Prox�y Sv��  V�LOAאigh-wSpe��Skiݤ/ ef.>�Hf�ٰ�mmunic��o{ns�
!
���urE�'�7�rt �F4�a�con�nect 2;�I�ncr`�stru����� SpK�AREL Cmd�. L��ua��O�AD*�=�Run-;TiưEnv� �yD;�(�el +��]s��S/W�.{��Licens�e����
����og�Book(Sys�tem)蔭�J�MACROs,~��/OffseS��Z�MHٰp��� j;73ΰMMR���l�35.f��ec_hStop��t��R� ize*�MiL��O� 2�7�x���0����miz��o}dM�witch�h���a�.�� v�ދ�Optm��49����fil��O�RD��0�g�� 8�496�ulti-�T������CPCM fun,�^�.sv�oO�Ğ�� �^�5�ReKgi��r��	�!2��ri��F�  H�59k�1�Num �Sel*�  74� H��İ Adjyu���adin���O� ,[���tat	ub��\У��������RDM Rob�ot��scovej� �d em(�:ٱn� SW��Servoٰs�����SNPX b���1��g P�Li�br���1ăڐ 9� ɰ.3�0g o��tE�ss�ag� f�"�@ e����"g���/I_�
�I�TM�ILIB���� P Firmn���^�F�Acc����0���TPTX���5w10.� eln����������H57�3�rquM�imgula��� 2�7Touz�PaxѩE1� T��6���&���ev.��IU�SB po����i�P�a�� 0\s�y nexcep�t��3 <� \h5�1 ����odu�V#��9��Q�VxN�k"6PCVL{&��^}$SP CS�UI�d���+XC���auҠWeb Pl���t? �#S ��\"	2�������S��&ު�V?8Gri=dplay��&�� ��8�-iRb".�� @ � R-20�00iC/165�¦ d+�+�lar�m Cause/�1 ed�<0:�As�cii����Loaqd��V4�3Upl�0�_CycL�c�m��ori����FRA�[�am�) tdt���NRTLi�3O}nݐe Helݨo 542*�PC`��4�`�]�1tr�ߵ48��ROS Ethv�t[����10\ҠiR}$2�D PkߵDER0>1�E����of�A��,ΰ�FIm��F�� �z��64MB D�RAMު�@:�9RF�ROA[�Cell03� ����shrQ
�B�Zc���ÍUk�p�� pide�Wty2L�s��|0\z�!C�tdѰ�.��@"Emai��li���+С\�� R0�qZ$GgigE�N�4OL�@Sup"��b�W3oa�~�cro�������4��QM��Fau�est�A>�j�� myiH9.dVirt��0W��0{&ImM�+T����}$Ko�l B�ui��n�յ'AP�L�&��MyV6� "\�0�*CGP�l��փ{RG�'p�{SB�UW�RQ�)K�&c�m\:��z��fX�)Oؒvõ(TA�&sp	oҠ-�B�&��
 I�f\E P�+�CB'f�g-��&" 5 �E��sv�b��Hvv�3��S_k��TO;�-�EH�f6.
�EN�vfx_z�)�V���tr>�)�hZ%.�F��& � ��r���*�G��&���њr����Hx��РJzCTIAc�pw4�LN�1�Mr�" #[��g�"��M�-�P2�~Tp�@����vxui�-�S�&�S�&�*4��W��2.pc�)V�GF��fxwʪV{P2AU \fx����N�if�u���"�in��VPB����)��s�D��*��a<s�F�5 M��s�I��c��{&Traİ��U~,p  ��<��2���RDp	�N���HY���p��-���H���Øp)����� �ϭ����yħ���rд��Ϟ�í4+���'�9L���ӎ��yy�9ӫ�c3ߞU��B�O�q�u���kߍӍSyy*�ߩ�\Yy�ߞ��k�W���ӄ��Yx����:�y	�������5�o�e/�Q���,�K�m��yg��^~��Ε�u�2��A��y������F������y�)���|�����1�m�.�<+�M��8G�i��7n��c���1�� ����W<�����7�{�����6�Z�������uk��[�|��!��?�ϔ��i�B\����_���{�x@.��wrst���B��� H68��@H�)T@J�EEND9I?��tql[}�
_�w�P�T�Q (��I) "���PA���T��/��85/A#b s;/�C/U/�,q�/�B�Gp�/�#��/�"3�6�5�R ?!2epai?5!:/Y4W���%INTo?e?_.�q�?4)��?�2pas2g�?�F O�?fA�ad6?��t Z�UD2gunOOqC5#33R?�D�0u�O�/��Mcm���OO�LNT�?��P_�Ĕ�0_0QR7�L_�Cfi._H?8_,_f'R50�_�S�AF-F�_�7�w.vo��_�_8�/�dM Cbo���o�bvrEo��paa��oaD�@�osF-A�S-sS�p'Is(8�PCesXPL�O�tslo_�ut\a�O�h%afvh%- B ��/����C�$��srp�?@_�?`w�"}�bA�����h�`���]T�ˏ�sgch��os�t��CG\s�;��us�?���Sg��/�G J����G�Dǟi$"�o�gdiʏ!�fd���?�h%J64S��Tut �o�O�?s����F�_夀���E�0���D`!��)�NO4E�O�i$II���iwjOl�ž0��>�?*�lb
��V��vjr/��
���7���ϥ�_�?zG7\ 2O�EG��Ϲ?���1՘ ޯ��_d�oi�8 ��c�50�>�x�Ͻ�"Lo�h%����dj9�﴿ƿؿ�c�� up9�C� j9�{�E��L��Ek, B串����oS_e_�&p/��O}�j94J���duZ��U��=d`;�����8���r7�Dhu���;]m T��������f�a���M���0�P�-4r V���O" #S�dwcL�P�in�`�a�?f& HTuRef�&��
�?hc�g�qr"��q.JG"�erM/��/ �/LsRA^��uH71�/��tCK�/<eTXP�/?i�k1/m5k.f���riR�eHG�/�/ cr�N'HGRf?L�iY�7�2hOuX��H\mO�� oρ�;H��DD@�O�� *�<�:I�?�?��d�R�η_ hd�ghg`OO�_���gmh�_h�m��XO�o|O�O�o��O\/�o0�f�gm �o`��`e۠;i�ov��yt��"��uRc60���#tmo�_�#1��fd r,op7��_�����lp>oh��冬'~ ߏ�dgts���&dޏ�/�o0�o
�J?<�vrF���cv.R���Ɵpld�56�%4�0/���greeK�m�XP)�fKCO*O|%56?��OZ� o~����E$i�o����jߠ���l ̂���OR��LOFvod��_IF��$��� ߪ�DߦX!B� Uc�e��t�4 ���(	M�O�5)e?Ƕ/���`1?Q�D�uk� '�|����`�boto�����-���6�p�eS ��on*���^� lB'����Տ_�q�_�rdk��4f��C( ҿȿ¯ԯ������̟p�����
I���571��t�ad�i39Tar��l�o�fk�������vPå@� PJ��|*���������e�t�4epg���ed��� E�5�RI�  H5�52� 747�2�1�pWelRK78�,� �0E�TXJ614���ATUP � wmfh 54�5�p�"6�pk��VCAM  7�\awCRI�@ ED" G UI�F)!28  j�CNREM�`��63�a�SCH�  4C DOsCV� CSUi��!0 D sEgIOCE�54�n#R694 we!!ESET=S#!3!�a� 73!fanu�MASK��OPRXY�_"7� ��0�OCO��"3�=P[�#"�ER J��" 7�!!J77�4#!39�  Eq8�G1�LCH 0#�OPLG%J50�00#MHCR)%P�S�17#MCS 4pD"�04 O#J55 �[#MDSWe!Y1M�D#1s#OP#1#MPR$07�0w"0�#8�  �#PCMX �#R0A�#� &�00��#� ( �&0�$50�( �#PRS� 3Js6903FRD@ �02RMCNy�n�dM�93 �SNBAA�80�0�@HLB  "�Lo�SM�A0 �(Ww"4 onitz#!2  II)��TC [#TMILpe �B�`0"K3�@�TPA� �QTXna�t\j�@EL�B&M250`0/D8��$�78�mon�19�5d SD95\FUEqC 0OP� UFR@ ���;!C@ \�@;!O:�0pt"VIP�@#� I�@0�!CSX�� �#WEB �#H�TT \stB2�4 �#CG�Q#IGޫQtopm�PPG�S!��PRC�@SH�7���w!6( �8���![�R RBB- sCi�B01rogw!f#IF#"098-!�!` �@�A64�(AaNVD�!Ld�1h 6a68( c�`d S{R7c!te.p� �0kaч@�bc`� CCLI$0?�sb$c9G �MS�"5a�` - �A� STY�@al� �@CTO �CJ�NN0J98�O�RS�0G��b�g �J�`OL�1Abn�: SENDu�to��!L�Q���@*r#S�LM� 8�"FVRn� MCHN0CSW!�SPBVP�� P%L� ds �qV$0�c�CCG $p�aCR҄0
Np�QB� 87�.f�QK� j70�*`�p�0'3CSqToo�CTQ���q�TB�P�N��@n$;pqC�@�Q#�� �p,#�p ��. %�$0h7#%� `8D#TC� QSQ"TE� [#m�, �tTE� gt"m�P�TTF�Q[����@�#CTG�Q�"���@ί#CTH `�TTI�@#CT'Qeqs�PCTM�@SC�$0xgS��0bodyq=P�@  ��� O�1� d��q�aus�a9��P[��qW `@06; GF� `8�V@VP2@ 6#23R i��@j?�g�R `n�g�B `" �g�D `��g�FX m;na"PVPI��+ �G V�!#V	`  23�RVK�@Np�@�CV�Q31�93{4.�vo R�erne땗�����i��r���h����A���37� ��"�\srv�����b�3b�- Sr�B"0���A�J935땿B�/5 (S�O���g �1�1�R|��j93땷b��ENz�5�� awm�{SK� Lib� �������� ���	 �"|�h�h��#��b�wmsk"�nE����q����pyE�  ���!x�02�t Fuï�բ6ۯm��uji%-�I&���8k�� 8!�Ń�땼P��2�p2�2�Mai'�on��_�/r�;pڦh;�;�G��_r���!v��4\ֶORC�ֺ+�5�� "T¦T�P��hQ�652�10��4���<�xk������ߦ�t�P��QrxֶSB�� ch_�����)�t!0�B�"̿ h�h땇�;���c��� ���������>�Rp� \toֶ3���#cl�W��2p�"� ���������F� ���b� Qt�a�϶0�t��ܐFsȒ�76t�p�t	� Ad����582��ob�|g*{�\a���FMQ ���A�mi1gֶ�I�or�w�I�j�rfm��F�c���@1�EYE&~� w���R����4�K2Х70.�E�ld,�C�� 1PTP]���..�"AD.�F�&83 k���ask���"�`4���۳dֶےv��ER~�7 R�ƀ�/�T�?)�e�rv�G?Y?k?}?�?�?ӹapa��	d��h��r�4�M��te��"��79!J�d/���G�p�ac�T��<�6�b�/� QO��$v�c>�,@Vg����e�YW��5/� BJ�h���R5:�d��Ɓ0�@��I_�raaj��e��he}ǔ$`��5(Xa�@��eqt榻�1Otdj��h,�_h�\	UI�/k�jo�FO��`^���aF��r��qW65q���K �'6ڦus W'�b,'��'?��n��MFR��;]�blf�ǯ�fr>���w�p�/�,��_U[ǀ�мn�x'_i� {�����O���pJ���X[@�o�in7L��O�9�\^ �� R����+mi�2״h �j��҇- �f�nt >�MA� H�I  �H5529� (�Cߑ21��le�R78�c�ߒ0�AcaJ61�4���0ATUqP�����545�t�-fl�6yE=�V�CAM�tFLX�CRId���o�U�IFULX �2u8��mo�NREu'���63��WQ��SC�H��Cn�DOCV��gϠCSU1�cx�r�0$�;EwIOC%tx\c��#54�oQ��9T�;��ESET�Temo�?�S�/��7S�{�M�ASK��70��PGRXY�T�`��7�ú`�OߐOCOe�\B?�3�ô`>��0{��?��|�-��on G?�39!'ߑõ� H82LC�Hd��@IOP�LG�tCGM?�0x��GЎ�MHCR�Gbo�S�/1_�CS4�7cgm��50T���?�5$�[���MDS�WMf.�D�����O�P��X/2L_�PR��K�����{����883n�CM��0iA,��0�Ő`~�=5#�\h88��+�?�D���.?���4J��0D�3��o�S4�����9��,i�FRDd�/2E/���MCN5�H93��K�SNBA�U"�R��HLB��SM�՛ñ�T���J52��SaߐTC4�\�T?TMILe��Pt���A|�TPA�^��TPTX��5��'TEL�ԫ�0䴈P���8�˳���K�9�5����95��88�8��UECd�rt �UFRd�__��Cd�2e-�VCO4��VIP�;���I�TAX~�CSX8�����WEB4�����HTT4�ka��2^T�2M/So�G#��QIG��< .��IPGS=t\rxFO�RC��aߐ7��/a��6D�s@>�R7 #��!��Oq�Ҥ��P ��Ҷ;�A���KÑ�$��0 "��4����N�VD4���#�Adaep��8D���68��ƻ�R7���P��D0���a��o�bܠ. CLI��l\-C����CMS�'��4�d; "ްSTY�[�CTOT�tl��N9N����ORS4�;��1 ��ltiΰOLS�( E���0�T���EL��6�@���9@ ���LM4�HV fo�VR���CS��wshc>�PBV4�쫁/�PL�
APVust>�CCG�4��0nCR�4 �H5��B���K�H573���?�<���\cms�#�7st.~TB���(! ��7�C�ԓ�<?"�awsh?"���I0?"��3�TCpd�K�A 4�\sl"AEĤpP��� 4�C[��"Ԥ8c��"4�(��CTF��c��"�n��CTG�73m#YG�THd�h� ��I��K�CTC�5�9m�CTM�5M𔴻�Q0��re\g�P���12��0�4�����%S��1]3MCTWd�9[@�_�GFd�SE]�P2d�t+��2�ա �2nd�ell��PBd�I���1Dd��a�1Ftap VPILd���CV�!Vq�:�UA��CVK�ۣ�CV#�core L���H"�Hp!�HK"�Hatc�J�H��4�I� �IL0H �I�2�H��H+2�IL��Y4=�H���Ie\1a�I�2 Z93�I{ �H�@NZ+��H 1��K#48�Z<A�Ht{�I l �Z;"�O�Fs\!�H�k"�H{"@o�F[�PZo�Z���J��Tok�РH��H\��Il�Z���Z2=[ng-[gT�oo�I�p�j(�njr�obt_�Xbt.�JL� iur�o�I� �i�!��F��POz�ling�j��y���Y"r^zۢ�I�p��Geat^j�]��Z��_je�����_��lkҠHm,��H|��Z���A�I  �_�s  ���Gvhm�J�{�svnj���H49�\�J�@L�Ij74u9{P�Zt\jNj��@_"g.pjmc3al�0�fu�J��^zhm-��_bg���o��\ͫ �1�H! �j��;����MT "�(Cu�zk��bg�ft�JlpX���GgCT"���Gfc]��˝26\fߟ�9C26�l\� Ίup�>m��;�Mul?��Q��7\^�K���7`-[˝���_�61Nj748.� H- �H��@R_�L^ziPe0��K�Я�F8\}�}�`����Ћ� � Rk,�ticMoj+@Oo�Qxs-@�"�3�CS� j+}LB-[5 9HNj+� co~�L�d�z��f�k˝lb��jll����-˜�k�/�.���LЎ�kipJ/�on,�J\A��]8�SK"�� ��wuto�o B��X����kwm� �o��Htp�ʜ n}��#ex-�˝��x���%a^jlL�je�식	i��a��/���{rej�1�o,�Vor�zR�����e T�Z[��[lc�lN��߭�SOžG3ZD��to�{+BΠH643N�`�SG/o��sg�a�Utui��;`�J��`��;�ndm�ndi N�{/�/�/�/�/�/�/��/??/?A?�?��r�iΪ! -Kj95�0/�n �zk]8915n/�O�t �Z���wsg�K,�>��i;ag� SGJ����ogu���KO]Lstw>_@	J64�:1�s�{F O>ګ#cdݛ��`3_��Yr-��N74�y-��3��RINnzlly��(m^���L����sgc�zI" #p?
+�oߡ\tw/� ��0.�@�"���f�_ʯ[y�Kmm�K}dc�t^�t]�+�
PR�ZWCHK
k, �;;`y<p��lK����LN*R85j ̛@_jR ���ti�N�g WJhecdN�L�F����wlZw|*�dat��Λ�greN��o�  STD��r7LAN-G�Aoc�e�`���Q�7��R87�0�{��8 (P�ogge����!�58\�PAcTTs�� �t\�N�c "B�@V�<�1�patd���O���������{q�
��5�a�p[�m�\q㕻�7�\aw��@�a��p6�����<ϯ�gmon���d��0�B�m�;A���\ ö��K�I�MH{CR�51 H��B��g\o��@��R]Ǐ H54ۿm�<@E����;!�����om�m�;a��R�|�N㕬0F�C��W�P�)Ai6�� Fƫ�{��itx�#{ ��icaio����De6��eve����72 �R�@RƜPg��ad�l��nt��K�RBT�tOP�TN`772'�CTK"'�g�(䔠�)� "AZ'�;q'圻q'�tzn&�{ E�'�Ama��- M�u��ncInDPN�������O872��|�d��(��������#����masy��y "�M��o��䃲��et����\p1�����\ 2��f���lZ����lp���9���`��+ V��ail��?������䓢��zd�<�k`���73.f��ir�dg��- i��ep\ ����� S0j�021"�1W ��(��`�4�� (i��e,"� "���+���/core_�I��l`aF��AY��AB���@����H�����AB;IC��Par;�M�ai������<� ;c\�ITX>����  ����1���g Jclib��ShiW�4��� t994\�V�SSF��� tt\{j9�f "O�pw� t��$%ini�/��pٰ t�5G�&�,� t\vsR&x�Lx�%w� tamclS/+ref.�%#� t	j��%m�� t[A�&�4\z�/�,z_v��%A�%�a�%_ol�6��l% �%end��/<c?.?@?R5o�[?m>�6�/�dshf�/+trt�?<O<AE�'F  !�G��$%��5vi�6���6� J92�F3��%2'5 (�%�@e&�Px�%k�4O dnwzFb��T�&`�XEpn�&|g��? nw\n�?&�,nd�V��N;XnF� j���%se�V I/
&�q&фU�n�5r w�%/F� X�F�_�rclR&0\p,w/Y�90�Eo`/:"5Of "U//A+dprm�%g¨%�XCrsu/kmS�T_ L`�6/OŔpM�LO�j��`nO1|h�ODnon8�|YCwrpR/�lp���E<�Pe\ga��Krgas�o�k�b�f�v��4xtfL�?m$ra�o�la00�omk�_�TamN6+�p4�`'9K0.v�W�ې�%�@�Ft��XE �sV��ДJ737�%|*�%,P���hB "+��Kwcf�F& I����998�vtomzFut  vV�_	o;�YC���:#8\F&�Y/� 0��f��deb^V��$@�0zFؠ"��g����<9\�&��9�Wrl}  �su"�st�G`��X �f� U (�fagn�F PzFϜ�V�ia�TX����v�d��w��g��HzF- O�W CH� �$G723�F���E(Aπÿտ2蚽Wc��Ws�vF& S�W�JR64��_�RVo RV���ӊ��vt�M\�etF�XoN�o�Fr ��x���+�1T�F?zteR� J58�O�  34	Wglea,�%,�j�Dq\t"���zFwIta1lUT�A�VϜ�gw韗Ma�d�W�Oa���6d �M��e�FT��90� H�%NT��R6�9������ir\�ʆMIR��ӊen�ʆv���F|�3��ITCP��Ta0�p����(MM7G�eT�o �\tpʆI��YBbusJ׈�m��I�@zFȀ��F�����/:��W�'g, ��4`�R_(!sw�&s_YC6c7\JF��Tf_�����Dfw��W��4a3chg��a96_���� _���_rV�% 99YA��e��$FE�AT_ADD ?_	�����?  	�$YA //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o #5GYk}� �������� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿�������DEMO �N�   ��*� �2�_�V�h� �������������� %��.�[�R�d����� ������������! *WN`���� ����&S J\������ ��//"/O/F/X/ �/|/�/�/�/�/�/�/ ???K?B?T?�?x? �?�?�?�?�?�?OO OGO>OPO}OtO�O�O �O�O�O�O___C_ :_L_y_p_�_�_�_�_ �_�_	o oo?o6oHo uolo~o�o�o�o�o�o �o;2Dqh z������� 
�7�.�@�m�d�v��� ����ƏЏ����3� *�<�i�`�r������� ̟����/�&�8� e�\�n���������ȯ �����+�"�4�a�X� j���������Ŀ�� ��'��0�]�T�fϓ� �Ϝ϶���������#� �,�Y�P�bߏ߆ߘ� �߼���������(� U�L�^������ ��������$�Q�H� Z���~����������� �� MDV� z������ 
I@Rv� �����/// E/</N/{/r/�/�/�/ �/�/�/???A?8? J?w?n?�?�?�?�?�? �?O�?O=O4OFOsO jO|O�O�O�O�O�O_ �O_9_0_B_o_f_x_ �_�_�_�_�_�_�_o 5o,o>okoboto�o�o �o�o�o�o�o1( :g^p���� ��� �-�$�6�c� Z�l���������Ə� ���)� �2�_�V�h� ������������ %��.�[�R�d�~��� ����������!�� *�W�N�`�z������� ���޿���&�S� J�\�vπϭϤ϶��� ������"�O�F�X� r�|ߩߠ߲������� ���K�B�T�n�x� ������������ �G�>�P�j�t����� ��������C :Lfp���� ��	 ?6H bl������ /�/;/2/D/^/h/ �/�/�/�/�/�/?�/ 
?7?.?@?Z?d?�?�? �?�?�?�?�?�?O3O *O<OVO`O�O�O�O�O �O�O�O�O_/_&_8_ R_\_�_�_�_�_�_�_ �_�_�_+o"o4oNoXo �o|o�o�o�o�o�o�o �o'0JT�x �������#� �,�F�P�}�t����� ����������(� B�L�y�p��������� �ܟ���$�>�H� u�l�~��������د ��� �:�D�q�h� z�������ݿԿ�� 
��6�@�m�d�vϣ� �Ϭ���������� 2�<�i�`�rߟߖߨ� ���������.�8� e�\�n�������� ������*�4�a�X� j������������� ��&0]Tf� ������� ",YPb��� �����//(/ U/L/^/�/�/�/�/�/ �/�/�/ ??$?Q?H? Z?�?~?�?�?�?�?�? �?�?O OMODOVO�O zO�O�O�O�O�O�O�O __I_@_R__v_�_��_�_�_�_�_m  h$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ ����"�4�F�X�j� |�������Ŀֿ��� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�t߆ߘߪ� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: L^p����� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲���������>�  �� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZl~���� ���/ /2/D/V/ h/z/�/�/�/�/�/�/ �/
??.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo Xojo|o�o�o�o�o�o �o�o0BTf x������� ��,�>�P�b�t��� ������Ώ����� (�:�L�^�p������� ��ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ�������� �*�<�N�`�r߄ߖ߀�ߺ����������	�,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oi��$FEAT_D�EMOIN  Vd�D`�`,d_INDEX9kHa��,`ILECOM�P O����zaGb'ep`S�ETUP2 P�ze�b�  �N �amc_AP2�BCK 1Qzi  �)h�o�k%�o`}`A e�om�o� �� V�z�!��E�� i�{�
���.�ÏՏd� �������*�S��w� �����<�џ`���� ��+���O�a�🅯� ��8���߯n����'� 9�ȯ]�쯁���"��� F�ۿ�|�Ϡ�5�Ŀ B�k�����ϳ���T� ��x��߮�C���g� y�ߝ�,���P����� ����?�Q���u�� ���:���^������ )���M���Z������ 6�����l���%7 ��[��� �D@�h��i�`P�o� 2�`*.V1R`� *c�`����JPC�|�� FR6:�".�4/�TX`X/ j/�U/�,;`%/�/��*.FM�/�	���/<�/<?�+STMG?q?��]?�=+?�?�+H�?�?�7��?�?�?EO�*GIF OOyO�5eO"O4O�O�*JPG�O�O�5�O�O�OM_�JSW_�_� �Sn_+_%
Ja�vaScript�_�OCS�_o�6�_��_ %Casc�ading St�yle Shee�ts0o� 
ARGNAME.DT_o
��0\so1o�Q�d��o`o�`DISP*�o�o�0�o7�e)q�8�o
TPEIN�S.XMLg:�\{9�aCust�om Toolb�ar��iPASS�WORD.�F�RS:\�� %�Passwor�d Config @����������� r�����=�̏a�s� ���&���J�\�񟀟 ����K�ڟo����� ��4�ɯX������#� ��G�֯�}����0� ��׿f������1��� U��yϋ�ϯ�>��� b�t�	ߘ�-߼�&�c� �χ�߽߫�L���p� ���;���_��� � ��$��H����~�� ��7�I���m������ 2���V���z���!�� E��>{
�.� �d��/�S �w�<�` �/�+/�O/a/� �//�/�/J/�/n/? �/�/9?�/]?�/V?�? "?�?F?�?�?|?O�? 5OGO�?kO�?�OO0O �OTO�OxO�O_�OC_ �Og_y__�_,_�_�_ b_�_�_o�_�_Qo�_ uoono�o:o�o^o�o �o)�oM_�o� �6H�l�� �7��[����� � ��D�ُ�z����3� ԏi��������ß R��v�����A�П e�w����*���N�`����֦�$FILE�_DGBCK 1�Q������ ( ��)
SUMMAR�Y.DG����M�D:3�s���D�iag Summ�aryt���
CONSLOGi�L�^��������Console log�����	TPACCN��R�%:�wς�T�P Accoun�tinρ�FR�6:IPKDMPO.ZIP�ϯ�
����σ���Excep�tion ߱�_�MEMCHECKm��Կb����Mem�ory Data|��֦LN�)n�RIPE�\�n����%�� Pa?cket LϺ���$SA���STA�T�����ߋ� �%�Statuys��<�	FTP�����r�����mment TBD���� =�)ETHERNEU���B��S�����Ethe�rn(��figu�ra߇���DCSVRF���������� verif�y all٣M�(��DIFF�����/di�ff�PB���CH�GD1�x�c �FQ&��	�2�� 85�YGD3���'/ �N/��UPDATES�.m S/��FRS�:\k/�-��Up�dates Li�st�/��PSRB?WLD.CM�/����"�/�/�PS_ROBOWEL1���:GIG�ߊ?/��?��GigE ~��nostic*�~ܢN�>�)�1HADOW�?�?�?�5O��Shado�w Change���٤8+�2NOTI��O"O�O���Notificx��\O٥O�A�� _��2_կ?_h_���_ _�_�_Q_�_u_
oo �_@o�_dovoo�o)o �oMo�o�o�o�o< N�or��7� [���&��J�� W������3�ȏڏi� ����"�4�ÏX��|� �����A�֟e��� ��0���T�f������ ����O��s����� >�ͯb��o���'��� K��򿁿ϥ�:�L� ۿp����Ϧ�5���Y� ��}���$߳�H���l� ~�ߢ�1�����g��� �� �2���V���z�	� ���?���c���
��� .���R�d�����������$FILE_�� PR� �����������MDONLY �1Q���� 
� �)�@_VD�AEXTP.ZZ�Z��p�G�L6%�NO Back? file !��U3�M��7� ���G�&�J\ ����E�i �/�4/�X/�e/ �//�/A/�/�/w/? �/0?B?�/f?�/�?�? +?�?O?�?s?�?O�? >O�?bOtOO�O'O�O��O]O�O�O_(_��VISBCK����*.VD)_s_�@�FR:\BPION\DATA\^_�R�@Vision VDt�_�O �_�__o_Ao�_Ro woo�o*o�o�o`o�o �o�o�oO�os� @�8�\��� '��K�]������� 4�F�ۏj����̏5� ďY��j������B� ן�x����1���ҟ�g���MR2_GR�P 1R����C4  B�O�	� 
������E�ˀ ֯�r���OH�cEP]��O���#M��
�KA���?�&�r����:6:N=�R�9-�Z���A�  v���BH���C`}dC��=N��B�{��r����пὫ�@UUT��U����/Ϫ��>��>c���>rа=ȫ��>i�=����>����:���:��:/�:6)�:��~ ϗ�2ϔ��ϸ�������z�_CFG =S��T  �a��s߅�0[NO ^��
F0�� ���/\RM_CHKT_YP  ���O�h���������OM���_MIN��L�������X��SSuB7�T�� ��5�L�,�U�g����TP_DEF_O�W��L�����IR�COM�Ѝ��$G�ENOVRD_D�O��	��THR��� d��d��_E�NB�� ��RA�VC��U�UQ ��Υm�X��|��������� � �O�U��[��O�x���⾥8�:����
,.  C�������h/�v%�������\n�!�SMT'�\.����+�w�$HOS�TC7�1]K[[�Y� 	MM�MI�}�e���� /*��1/C/U/g/��/ 	�anonymou�s�/�/�/�/�/?  L^pM?�/� /�? �?�?�?/�?OO%O 7OZ?�/�/O�O�O�O �O? ?2?D?FO3_z? W_i_{_�_�_�?�_�_ �_�_o._dOvOSoeo wo�o�o�O�O_�oo N_+=Oa�_r �����o�8o� '�9�K�]��o�o�o�o �������#�5� |Y�k�}�����ď� ������1�x��� ��J��������ӯ� ��	���-�?�Q�c��� ��Ο����Ͽ��:� L�^�p�Mτ����ϕ� �Ϲ��������%� 7�Zϐ���ߑߣߵ� ��� �2�D�F�3�z� W�i�{��������� �����
�d�A�S�e��w����/ENT {1^�� P!�.��  ���� ��*��Nr5~ Y������ 8�\1�U� y�����4/� X//|/?/�/c/�/�/ �/�/�/?�/B??N? )?w?�?_?�?�?�?�? O�?,O�?ObO%O�O�IO�OmJQUIC�C0�O�O�O_�D1 _�O�OV_�D2W_3_�E_�_!ROUT�ER�_�_�_�_!�PCJOG�_�_�!192.16?8.0.10�O�C?CAMPRTGo#o�!7e1@`noUfR�T�_ro�o�o��NA�ME !��!�ROBO`o�oS_�CFG 1]��� �Au�to-start{ed��FTP��~q���F��� �����9�K�]�o� ���&���ɏۏ�����#���Wi{X� ���o�����ğ֟�� ����0�B�e��x� ��������ү������ �Q�>���b�t����� ��q�ο����9� ��L�^�pςϔϦ�� �����%��Y�6�H� Z�l�3ϐߢߴ����� ��}��� �2�D�V�h� ��������������� 
��.�@��d�v��� ������Q����� *<������� ��������8 J\n��%�� ���EWi{} O/��/�/�/�/�/� �/??0?B?e/�/x? �?�?�?�?�?/+/=/ �?Q?>O�/bOtO�O�O �Oq?�O�O�O_'O(_ �OL_^_p_�_�_(�`_ERR _z��_�VPDUSIZW  9P^S@��T�>�UWRD ?�EuA�  guest3V�$o6oHoZolo~o�dS�CD_GROUP� 3`E| Iq�?YM �nCON��nTAS�nL��nAXP�n_E�o9P�n��RTTP_AU�TH 1a�[ �<!iPendCan�g�~@}9PJ��!KAREL:q*���}KC�����pVISI?ON SET�`E��I�!\�J�t��s�� ��������Ώ��-����dtCTRL �b�]~�9Q
9QFFF9E39��DFRS:DE�FAULT���FANUC We�b Server ����dtodL��'��9�K�]�o��TWR_~�`FIG c�e��R���QI�DL_CPU_P5C9QB�@�w BHǥMINҬ��a�GNR_IO�Q�R9P�XɠNPT_SIM_DO��!�STAL_S7CRN� �y�+��TPMODNTOqLY�!���RTY8�p�&�9�hpENBY���cƣOLNK 1d�[�`������1�C�U�ͲMAS�TE���&�OSLAVE e�_|˴jqO_CFGs�Ʀ�UOD��Ϩ�CY�CLE�Ϧļ�_A�SG 1f���Q
 W�9�K�]�o߁� �ߥ߷����������8#�_��NUM�S�bz�U
��IPCH���j�O_RTRY_�CN��Z��U�_�UPD�S���U ������g�θ`����`ɠP_MEMB?ERS 2h��` $�e�>���HyɠSDT_IS�OLC  ����r�\J23_DS�q���OBPRsOC��%�JOG�d�1i��89Pd?8�?�.���".�?�?�?OQNs ��V����3W~����������POSRE��$�K_ANJI_m�K��i�pMON j�k~�9Ry���� //�^�r��k����a9%Th��p_L��I�l�kEYLOGWGIN���`�����U�$LANG?UAGE ������ �!�QLG���lq�9R��9Px^�p�  ��砭�9P'03X�k����MC:\RS?CH\00\��� �N_DISP �m��DAMK�SL�OCw�آDz ���A�#OGBOOKG n���9P~��1�1�0X�9O%O 7OIO[OmN�Mɱ���I��	�5Ib�5�O��O�5�2_BUFoF 1oؽ�O2A5!_�2��=_?7Y_ k_�_�_�_�_�_�_o �_o:o1oCoUogo�o��o�o�oe4��DCS� q�= =��͏L�O-�1CUg|���bIO 1r�G ��s20� �������1� A�S�e�y��������� я���	��+�=�Q�Z|uE�TMl�d ����Ο�����(� :�L�^�p����������ʯܯ� ���7�S�EV��u={�TYPl���z�����!��PRS���/S��F�L 1s�}��� �$�6�H�Z�l�~�F��TP� l�i��=NGNAM��A5�"ne4UPSm0GI���\!����_LOA�D��G %u:%�REQMENU���3�MAXUAL�RMI�c�W�T���_PR����3�R�Cp0t�9�M���3xEݗ���P 2u��W �1V	i�00���߭�1� �.�g�xU���� ����������8�J� -�n�Y���u������� ����"F1j M_������ �	B%7xc �������/ �/P/;/t/_/�/�/ �/�/�/�/�/�/(?? L?7?p?�?e?�?�?�? �?�? O�?$OOHOZO�=O~OiO�OK�D_L?DXDISA�����zsMEMO_AP���E ?��
 b��I�O_"_4_�F_X_j_|_R�ISCw 1v�� ��O �_ ���_�_�Ooo�@o�_C_MSTR� w:�_eSCD 1x�M�4o�o0o �o�o�o�oP ;t_����� ����:�%�^�I� ��m������܏Ǐ � �$��4�Z�E�~�i� ����Ɵ���՟� � �D�/�h�S���w��� ¯���ѯ
���.�� R�=�O���s�����п ����߿�*��N�9��r�]ϖρϺ�PoMK?CFG ynm��~��LTARM_��z�����и����6�>�s�METPUl�ӫІ�viND��ADCOLXի�c�oCMNTy� l�g` {nn��-�&������l�POSCFz����PRPM�߶��STw�1|�[� 4@�P<#�
 g��g�w��c��� �����������G� )�;�}�_�q������������l�SING_�CHK  |�$_MODAQ�}����W��#DEV }	�Z	MC:W�HSIZE�M�P��#TASK %��Z%$123456789 ��!TRIG 1~�]l�U%�\!�S
K.�S�YP�69�"EM_INF� 1� �`)AT&�FV0E0X�)��E0V1&A�3&B1&D2&�S0&C1S0=>�)ATZ�#/
$H'/O/�Cw/(A/�/b/�/�/�/? �&?���/�? 3/�?�/�?�?�/�?�? "O4OOXO??�OA? S?e?�O�?�?_CO0_ �O�?f_!_�_q_�_�_ sO�_�O�O�O�O>o�O bo�_so�oK_�owo�o �o�o�_�_L�_o #o��Yo��� �o$��H�/�l�~�1 ��Ugy���� � 2�i�V�	�z�5��������ԟPNITOR��G ?k   �	EXEC1T���2�3�4�Q5�� �7�8�9���������� (���4���@���L��� X���d���p���|���U2��2��2��2��U2��2Ũ2Ѩ2ݨU2�2��3��3���3(�#R_GRP�_SV 1��� (��  ��m��MO�_Ds�����PL_NAM�E !����!Defaul�t Person�ality (f�rom FD) ���RR2�� 1��L6(L?�<���	l d��n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲�����B2]�� �*�<�N�`�r�����<��������� �,�>�P�b�t������BJ  ��\  �  ���Ȱ�  A��  B��T���� 
��������  ������Bz��p���  CH �CH P Ez�  E�� E�/` E�;%Z�Z�*� ?�  E��F��@&��T
 Ai� dx� H�x�	$Hxd�dڭ�}` (d��8(xx$$y Xt$d D (DDd pWwX��	X��vXHX���/�y�y (� !0��  7%E	��Em�Xw$%XH$%P�� �/�/�/ �/�/�/??+?=?O?a?s=F�r?�?�?��?�6��E�{P�EU���2 ��B�����?Kزd��'O9NO\OjG�0���|M��'4 � W%�O�O�N  �H�O�J�A  A��C�����_�OC_9W�  � TB�LY�@
��_�\B�@Q�Y=�CÈ��V�`HR0� ʒP( @7%?��a�Q�?ذaر@�6��&س��2n;�	l�b	  ����pX���U�M`�X� � � �,� �rb�@K�l,�K���K��2�KI+�KG0�/K �U�L2o�E�	O�n�@@6@� t�@�X@�I��b`�o�C��N����
���}v������` q�m�|�kQ�
=ô��  Hq�o~`!b���  Ȱ�a� �B����ذa�s�G��}�m��o�q��v�O��E	'� � 0��I� �  �� Q�J:�È~T�È=���l� �@|���}~�Q����R ����yN8���  '�<�ap?���b!p��b){�B��?�C�IpB  X��ذ���C�A�f��՚n`��(��BB P��8�����P��ԕرD �O���O���A�,�>�Š
��`l�1�	 S٠p��� p` l`�:GT  �t�?�ff{O��įV� �P���=�a�!��/�?Y)R�a4�(ذ]�Pf����a\c\d^ƃ?333-d�<��;�x5;��0�;�i;�du;�t�<!�+}�oݯ��b�Sb�P�?fff?��?&���T@��A{#$�@�o[,� ��x�	�&f6�ed�g ���Hd㯸ϣ�����  ���$��H�Z�E�~���&eF��mߺ�i߀��U���y���2���E�0����y�d�� ������������ ?�*�܏r�8�.o�ߺ� ���T�);ڿ Pb��������P��A��T C�=�ϵ��Y}��2������m�C��W�C�= �` Ca��������(!�`�<����bC@_;C9��BA��Q�>V{È�����Y�?uü��
/�S���Q��hQ��A�B=�
�?h�Ä/iP�����W��ÈK��B/
=�����Ɗ=�K��=�J6XK��r#H�Y
H}���A�1�L��jLK����H:��H�K��/0	b�L �2J��8�H��H+UZBu�a?�/^? �?�?�?�?�?�?O�? O9O$O]OHO�OlO�O �O�O�O�O�O�O#__ G_2_k_V_{_�_�_�_ �_�_�_o�_1oo.o goRo�ovo�o�o�o�o �o	�o-Q<u `������� ��;�&�K�q�\���΀�Gϭ���� C�aɏ Ĉ�y���CVF������+b�����yKc�f�� 
E��Ў�T�ٟ��(���_3�h۟���������N�������3�lC�(�:�H�����T�f��t�.3礁}����k����q'�3�JJ �����گ���4�"�J]P̲Pf��������⟛�ſ���ԻA����/��?�{?�<N�u�  fUh�*� �Ϟ������Ϣ�t�.��R�@��X�bߘ�̆ߨ�)Z�ߺ�  ( 5�	�������B�0�f�t�  �2 E%p"E[[@��N�"B,C��%@ߏ����������3�E�c������@����%n�n�%�đ�%��Xc
 ��!3EWi {��������b*[��P�I��v�$MSKCFMAP  ��� ^������pDONREoL  X�[���DEXCFEN�B�
Y�FN�C��JOGOV�LIM�d��d�DKEY��%_PAN�""�DRUN�+S?FSPDTYw��<��SIGN���T1MOT���D_CE_GRP� 1���[\ ���/��?&?��?Q? ?u?,?j?�?b?�?�? �?O�?)O;O�?_OO �O�OLO�OpO�O�O�O _%__I_ _m__f_��_O�DQZ_ED�IT�$UTCO�M_CFG 1�BQ�_o"o
�Q__ARC_�X���T_MN_MO�D���$�UA�P_CPLFo�N�OCHECK ?=Q W��� �o�o�o�o'9 K]o������vNO_WAITc_L�'�W� NT�Q��Q���_E�RR�!2�Q���� �_t��������*��Ώ�d``OI���P�x ���_ � ´ӏ8��?0�4����d�B�P�ARAMJ��Q��������s��� =��345678901��� � ��?�Q�-�]�����u�0��ϯ����������7�ODRDS�PEc�&�OFFS?ET_CAR�PKo�m�DISz�K�PE?N_FILE���!�$a�V<`OPTIO�N_IO
/!аM_PRG %Q�%$*	�ά�WO_RK ��'�� ��K�7U��h��f�(�f�	 a���f�7���M��RG_DSBL  Q�����L�RIENTTO* ���C�Y��M�UT_SIM_Dط�X+M�VQ�LCT �%��R_�$a<Q�'�_PEXh`��nb�RAThg d��b�r�UP �5� � ����߼߬����$��2�#��L6(L?�>�	l d'�O� a�s��������� ����'�9�K�]�o� ��������H�2>��� ��/ASew�N�<������ �1CUgyjH���P�� ��  ��  ��U�A�  Bl��PB����}H��  ���VU�B�p�������N�P Ez�  E�� E�/` E��;(�Z���Z�/��?�  E��''����@#���T
�AJ(��E!Y!a! )!m!Y!u)%)!Y!E!�%E!ڎ$�^$A!� 	!E!a!�%%	-Y!Y%�-58�Z 99U%$E!�D!	$D%%E! Q481X291�%�)95�/�W#95)%91m5a!�5/�Z7��Z (�8�10�<a1 EE	�(�Em�494X6E9=)%E15�� |O�O�O �O�O�O�O�O__0_B_T]F�S_y_�_�_�Vh�����_�[��%�on�_=oKg��]�]&�'4 ?� W%po�o�X� g��g�o�jA��A��c����P�o�o$w���tB�(~�`��r�|��� q�y�$�O��1��k����3�`��0���P(C @ED�D��q?Q��C�Z7}��o  ;��	lD�	u� ����p�X�[�2���X � � ��, �W��`H���9H�H����H`�H^yH�R�l���_h�����`C#�B�� C4ӄ�������9���
=��� ������c�Bz��Βa�m�另b��s�� �q���g䟒����Ǒ�ٖ�o����	'� � ��I� �  ��q<�=���89�K���@a�g� b���������唠�䮟�N��  '۰��Ɓ"�B�Ղ���т6��� �  ϥ�C�a�������`��2g�Bp��Н����px����D��o޿�o`��&��o�5���`Q��	 �٠U�f� U� �Q�:���#����?�ff\o�ϩ�;�C �p����"�8� ,��?Y
r��q=�	(� B�PK�fɆ�A��A���?333���m�;�x5;���0;�i;�d�u;�t�<!�!�y������t���r��p?fff?x�?�&��j�@��A�#	�@�o[ �	]����g��uI� �wh���-��ϝ���� ������	���-�?�*� c�u�L�������4�V�X��B�EjP f��^I�m� ��� �$�� W�������9 ��/ /��5/G/� z/e/�/�/�/�/�`�cA��$�t�/ C�/�"?i��Հ>�?�@�Pn?�/�?}?��(���W�?C�@�`C CT��?�j4�j0�i1A@I�!����bC@_;C9��BA��Q�>V`.È�����Y�?uü��
�?k����Q��hQ��A�B=�
�?h��iOJp�����W��ÈK��B/
=�����Ɗ=�=K��=�J6XK��r#H�Y
H}���A�1�=L��jLK����H:��H�K��O�@	b�L �2J��8�H��H+UZBu�?F_�OC_ |_g_�_�_�_�_�_�_ �_o	oBo-ofoQo�o uo�o�o�o�o�o�o ,P;`�q� �������� L�7�p�[�������� ȏ�ُ���6�!�Z� E�~�i�{�����؟ß ��� ��0�V�A�z��]9Gϭ���� C�a�/�� Ĉ�y�ЯׯCVF������üKG�j���yKH�K�� 
Ep��s�9���90(91�_3�h��y����i���N����LA3�lC���-¢���9�Kϰt�.3礁}e�w�k����q'�3�JJ �͑��Ͽ�������JB5P��PK�Zg�t�ǿ�ߪߕ��߹�A��������$�{$�<3�Z�  fUM�� ��������Y��7�%��=�G�}��k���)Z����  ( 5�� �������'KY  �2 E%pIFE[[@tN�IFB�!,�!� C��0� L@@į����*H3��Tfx���LCLB94���L@D=4H;
 �//*/</N/`/ r/�/�/�/�/�/�/�/�GJ@2��5�I��v�$PARAM�_MENU ?���� � DEFP�ULS��	WAITTMOUTT;�RCVg? �SHELL_WR�K.$CUR_S�TYL���<OsPT��?PTB�?��2C�?R_DECSN_0<�L	OO-O VOQOcOuO�O�O�O�O��O�O�O_._)1SS�REL_ID  ���Y�=UUSE�_PROG %�8:%*_�_>SCCR�k0ORY@3�W_HO�ST !8:!�T�_�ZT\Ю_ c�_��Qc<o�[_TI�MEi2OV�U)0GDEBUGMP8;>S�GINP_FLM1S`�gn�hTR�o�gWPGA�` �lC��kCH�o�hTYPE5<A)_#_Y �}������ ���1�Z�U�g�y� ������������	� 2�-�?�Q�z�u��������ϟ�
��eWO�RD ?	8;
 �	PR�`���MAI@��SU��1E�TE#`���	9�4R�COL��n����vTRACEC�TL 1���.B1 I�W֯|ࢵ�DT Q�����РD � ;��*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>� P�b�t����������� ����(:L^ p�������  $6@�bt �������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n�V� ������"�4� F�X�j�|�������ď ֏�����0�B�T� f�x���������ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰��ߘ ����
��.�@�R�d� v����������� ��*�<�N�`�r��� ������������ &8J\n��� �����"4 FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?�?O�C�$PGTRA�CELEN  �A  ���@�$F_UP ����SA�[@?A  T@$A_�CFG �SE�=CAT@��D��D�O�G6@�OhBDEFSPD �sL�A6@�$@H_�CONFIG ��SE;C @j@dT�3B A�QP�D�A1Q@��$@INk@TRL ��sM�A8�EFQP�E�E�W�pSA�DQ�ILIDlC��sM	�TGRP �1�Y l�AC%  ��l��AA��;H�{N��R���A!P�D	� a3C	\�T�Ai)iQP� 	 �O4VGgCoG ´|c^oGkB` �a�opo�o�o�o�o�b"�Bz�o�7I~3 <}�<�oN�J� ����f�)��9�_�J�`z����@
t���d�ŏ�֏� ��3��W�B�{�f�x�@����՟�����J)@�)
V7.10�beta1�F �@�@ㅟA&ff�Q2�C�PC�`�D�Dk�`[�C�T��@ �DĠ Dr� ��QBH�`�L��PC�5R A?�  F��CCx����b��P`!P��A����Ap`B��bc ��$�6��eC�QKNOW_�M  �E{F�TSoV �Z(R �C������ʿ��ٿ��$�A!m�SM�S��[ �B�	�E���Ϗ��*�E`��2�E@�2���������d@�QMR*�S�Y�T�j���A�Cf���e@�Rۚ]S�T�Q1 1�SK
 4�U��,ժ߲C �ߡ߳���������-� �1�v�U�g���� ���������	�N�-�(?�Q�p�2{���AG�<�����P3��������p�4��+p�5HZl~p�A6����p�7� $p�8ASe�wp�MAD0F �[E��OVLD  �SK�ϼOr�PARNUM  /|]///T_SCH� [E
}'F!�)=C�%UPDF/X%5U�/��_CMP_O�0@T@�@'{E�$ER_CHK5yH!6
?�;RS�]��Q_M�O�o?�5_k?��__RES_GzФ~� ���?�OO�?%OO*O [ONOOrO�O�O�O�O@�O�O��3���<�? _�5��(_G_L_�3G  g_�_�_�3� �_�_�_ �3� �_o	o�3@$o CoHo�3�co�o�o�2�V 1�~կ1e��@c?��2THR_INR�0�!7³5�d�fMASS �ZwMN5sMO�N_QUEUE C�~�f��0���4N0UH1NEv6;�p�END�q�?�yEX1E��u� BE�p�>�sOPTIO�w�;��pPROGRAM7 %hz%�p�o�l/�rTASK_I���~OCFG �hZ/\���DATuARè��@��2�����#�5�G�� k�}�������^�ן�x�����INFOR��܍�wtȟe�w��� ������ѯ����� +�=�O�a�s�������л�Ϳ(�4��܌ ��I��� K_���8��T��ENB� ͠�1>ƽ�I��G��2��� P(O8�ҡϳ� ������_EDIT ᭘��ߋ�WER�FL�x�cm�RGA�DJ �8�A�  h�?�0t�
qL��q���5��?�!��<@�x"*�%���@�#ߊ�f�2���F�	Hp�l�G�b��>�㻎A�d�t$I��*X�/Z� **:c�0V�h���Ǟ���B�����x"��� ����������b�� �L�B�T���x����� ����:����$, �Pb���� ���~(:h ^p������ V/ //@/6/H/�/l/ ~/�/�/�/.?�/�/? ? ?�?D?V?�?z?�? O�?�?�?�?�?rOO .O\OROdO�O�O�O�O �O�OJ_�O_4_*_<_ �_`_r_�_�_�_"o�_ �_ooo�f	���o �p�o�o�dJ��oL��o�#�oGY��PREOF ����p�p�
L�IORITY�����P�MPDS1P�>ߴwUTz�4�K�ODUCTw�e8�\�OG찇_TG;�|����rTOENT 1���� (!AF_�INE�pp�{�!�tcp{���!�ud��ˎ!�icm�����rXYڏӴ����q)�a p�/�A��p�)� j�M�Y���}������� �ן���8�J�1�n�HU�����*�s�Ӷ}}������,�>�%�
jfp�/z�֯K�,�������A��,  �p�������ʿ�u"�ut�}�sF��P�PORT_NUUM�s�p�P��_CARTREP��p��|�SKSTAv�w K�LGSm���������pU�nothing�Ͽ������c{t�TEMP ����ke���_a_seiban0C�,S�y� dߝ߈��߬�����	� ���?�*�c�N��r� �����������)� �M�8�q�\�n����� ����������#I 4mX�|�������3��VE�RSI�p �d �disabl�ed>SAVE ���	260_0H721:&��!;���̏� !	(�rmoN+E/`Áeb/�/�/�/�/�*�z,�? %`���_�-� 1����E0�b8eO?a?4gnpURGE_ENB3���v�u�WF�0DO�v��vWi��4�q*��WRUP_DEL�AY �CΡ5R_HOT %�f��q:�.O�5R_NORMALH
�OrOAGSEMIQOwO�O�lqQSKIP-3���>3x$�O _1_ C_]&ot_b_�_�_�_ �_�_�_�_o(o:o o ^oLo�o�o�olo�o�o �o $�oH6X ~��h���� ���D�2�h�z������$RBTIF��4G�RCVTMO�U\�����D�CR-3��I {�Q/ Qʴ1�Ed��A]	�C���3=;4~_  �j��QU�����_e�P�;��x5;��0;��i;�du;�t�<!��h��R���̝���� �&�8�J�\�n�����������RDIO_TYPE  4=���¯EFPOS1w 1�C�
 x/ :�H2��b�M���/�� E�οi�˿ϟ�(�ÿ L��pς��/�i��� ���ω�߭�6���3� l�ߐ�+ߴ�O����� �ߗ���2��V���z� ��9����o���� ���@�R�����9���������OS2 1��;+�u���-��xQ���3 1������G���gS4 1�~����ZE~�S5 1�%7q��/>�S6 1Ũ���/�/o/�/&/S7 1�=/O/a/�/?�?=?�/S8 1� �/�/�/0?�?�?�?P?�SMASK 1��߯ )�OF�7XN�OܯFUO_C�M�OTE���X4uA_?CFG �|M�1�\A�PL_RAN�GxA���AOWER� ���@�FS�M_DRYPRG %�%y?!_�ETART ��N�/ZUME_PRO��O_�_X4_EXE�C_ENB  <����GSPDdP�P8�X���VTDB�_�Z�RM�_�XIA_O�PTIONφ�����pAINGVERmS.a�z_��)I_AIRPU�R�@ @O�o�=MKT_�0T�@zO���OBOT_ISO�LC=N�F�1�a^�eNAMERl�bo��:OB_ORD_�NUM ?�H��aH721w  V1wLqrǈqrV0qr�sps�u\@��P?C_TIMĖ���x��S232�B1�����aLTE�ACH PENDcAN΀�7\H���x?c�Maint�enance C�onsV2�#�"��_�No Use��N��r�������8��С�rNPO>P�r�\A<e�qCH_�LgP�|Nw�	�<��!UD1:�b�	�R�0VAIL�Rq2e��upASRW  �:a�B��R_INTVAL1f��I�+n���V_DATA_GRP 2���qs0DҐP�?`��?�� o��������կï�� ���-�/�A�w�e� ���������ѿ�� �=�+�a�Oυ�sϕ� �ϩ��������'�� K�9�[߁�oߥߓ��� �����������G�5� k�Y��}������� �����1��U�C�e� g�y��������������	+Q?uDA��$SAF_DO_PULS�pE@�C��� CAN�r1f��vpSC�@���Ƙ�Q�V0D��D�qL�L�+AV2  y�'9K]o��������ڈ���2($Md�($C!u�1#
) @�Co/�/�/�.W)k/� M��$�_ @݃T:`�/??�&?39T D�� 3?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO�jO|O֏��i%�O�O�O܉�!L� ��;�o݄�p��M
�t��D�ipp�L��J� � ��jL���j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:����/c�u������� ��Ϗ��B�%�1� C�U�g�y���������Ƒ��0RMS�EW] �$�6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ��M���*�<�N�`� r߄ߖߨ�������� ��&�8�J�\�ǟ�� �������������� ��,�>�P�b�p��� ������������ %7I[m�� �����!30EWit�OB3 t�����// //A/S/e/w/�/�/�/�/�/�*��/?6���\R?�M	�1234567�8XRh!B�!̺��� �?�?�?�?�?�?�? OOA�>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_o]-O�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�oq_BH�o�o�o !3EWi{���������v[;�j�A�S�e�w� ��������я������+�=�O�a�xYD� k�������ɟ۟��� �#�5�G�Y�k�}��� ����v_ׯ����� 1�C�U�g�y������� ��ӿ���	�ȯ-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� σߕߧ߹������� ��%�7�I�[�m������v6�����z��!�3�O:C�z  A�z  W �@�2�v0�� @�
���  	�r������X������ph�u�����K]o�� ������# 5GYk}��0 ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-?G��������*@  <X4t���$SCR_GRP� 1�� ��� t ��t� E5	 �1��2�2�4��W1G3�;�97�7�?�?OC���|�BD�` D���3NGK)�R-2000iC�/165F 56/7890��E��?RC65 �@�?
1234�E�6�t�A�����C �1F�1�3�1)�1A�:�1�I	��?_Q_�c_u_�_���#H��0 T�7�2�_��?�_�_o�6�t���_Lo�_poB8boK�h��@��9BǙ�B��  B�33BAƿ`�e�b�c�1Ag���o  @t��e�1@<>@	  ?�w�b�H�`2�j�1F@ F�`\rd[o� s������� *��k�c)rU�@�R�d�v�B����ʏ��� ُ����H�3�l�W� ��{���Ě2C�?���7���9�t�!q=@"p6��G?�S��r�`y��`ȏ�@�G�L�3��ϯ�A>G��1��"oe��)�t� �<�N�\�*��q�}���^� P���(����ӿ�g1E�L_DEFAUL�T  �D���t���HO�TSTR� ��M�IPOWERFL�  K����?�W�FDO� S�R�VENT 1�����P0� L!�DUM_EIP�翬��j!AF�_INE��ϵ!'FT�������9!�_B� ��i��!RPC_MAINj�LغXߵ�|�'VIS��Kٻ���o!TP��PU����d��M�!
PM�ON_PROXYN��e<���g���f����!RDMO_SRV���g��1�!R�DM���h, �}�!
~�M����il���!RLScYN�@����8��>!ROS��<��4a!
CE>�MTCOMb���kP�!	vCO�NS���l��!}vWASRC ����m�E!vUSBF��n4�0� �����/�'/��K//o/�RVI�CE_KL ?%��� (%SVCPRG1v/�*�%2�/�/� 3�/�/� 4??� 56?;?� 6^?c?� 7�?�?� H�D�?�,9�?�;�$ H�O�!�/+O�!�/SO �! ?{O�!(?�O�!P? �O�!x?�O�!�?_�! �?C_�!�?k_�!O�_ �!AO�_�!iO�_�!�O o�!�O3o�!�O[o�! 	_�o�!1_�o�!Y_�o �!�_�o�!�_{/�"�  �/� F�E1��� �����
�C�U� @�y�d���������� Џ����?�*�c�N� ��r��������̟� �)��M�8�_���n� ����˯���گ�%� �I�4�m�X���|������ǿ�ֿρ*_D�EV ���oMC:�H'�?GRP 2ׇ�+p�� bx 	�/ 
 ,y�ϒ� +r~ϻϢ�������� ��9� �]�o�Vߓ�z� ���߰������#�z� G���k�}�d����� ����������U� <�y�`���������*� ��	��-QcJ �n����� �;"_FX� �������/� /I/0/m/T/�/�/�/ �/�/�/�/�/!??E? W?�{?2?�?�?�?�? �?�?O�?/OOSO:O LO�OpO�O�O�O�O�O _^?�O=_�Oa_H_�_ �_~_�_�_�_�_�_o �_9oKo2oooVo�ozo �o�o _�o�o�o#
 G.@}d��� �����1��U� <�y����o��f�ӏ� ̏	���-�?�&�c�J� ��n��������ȟ� ���;���0�q�(��� |���˯���֯�%� �I�0�m��f������ǿ������#�d ��	�4��X�C�|�gϠϯ�%����������������� ���+��O�=�s߁� �Ϧ���i��������� �	��Q��x��A� �����������Y� �P���)���q����� ������1�U���I ��Ym���	 �-�!E3U {i����� �//A///Q/w/� �/�g/�/�/�/�/? ?=?/d?v?-?O?)? �?�?�?�?�?OW?<O {?OoO]OO�O�O�O �O�O/O_SO�OG_5_ k_Y_{_}_�_�__�_ +_�_ooCo1ogoUo wo�_�_�oo�o�o�o 	?-c�o��o S�O����� ;�}b��+������� ��ɏ�ݏ�U�:�y� �m�[��������ş �-��Q�۟E�3�i� W���{����دꯡ� ï���A�/�e�S��� ˯���y��ѿ��� �=�+�aϣ���ǿQ� �ϩ����������9� {�`ߟ�)ߓ߁߷ߥ� ������A�g�8�w�� k�Y��}������ ��=���1���A�g�U� ��y����������	 ��-=cQ��� ���w���) 9_���O� ���/�%/gL/ ^//7///�/�/�/ �/�/?/$?c/�/W?E? g?i?{?�?�?�??�? ;?�?/OOSOAOcOeO wO�O�?�OO�O_�O +__O_=___�O�O�_ �O�_�_�_o�_'oo Ko�_ro�_;o�o7o�o �o�o�o�o#eoJ�o }k����� �="�a�U�C�y� g�������ӏ���9� Ï-��Q�?�u�c��� ۏ��ҟ�������)� �M�;�q�����ןa� ˯��ۯݯ�%��I� ��p���9�����ǿ�� ׿ٿ�!�c�Hχ�� {�iϟύ��ϱ���)� O� �_���S�A�w�e� �߉߿����%߯�� ��)�O�=�s�a���� ���߇�������%� K�9�o������_��� ��������!G�� n��7����� �O4F�� g�����'/ K�?/-/O/Q/c/�/ �/�/��/#/�/?? ;?)?K?M?_?�?�/�? �/�?�?�?OO7O%O GO�?�?�O�?mO�O�O �O�O_�O3_uOZ_�O #_�__�_�_�_�_�_ oM_2oq_�_eoSo�o wo�o�o�o�o%o
Io �o=+aO�s� ��o�!���9� '�]�K��������q� ��m�ۏ���5�#�Y� ������I�����ßş ן���1�s�X���!� ��y���������ӯ	� K�0�o���c�Q���u� �������7��G�� ;�)�_�Mσ�qϧ�� ��ϗ�ߓ��7�%� [�I���Ϧ���o��� �������3�!�W�� ~��G��������� ��	�/�q�V������ w�����������7� .����O�s� ���3�' 79K�o��� ���#//3/5/ G/}/��/�m/�/�/ �/�/??/?�/�/|? �/U?�?�?�?�?�?�? O]?BO�?OuOO�O �O�O�O�O�O5O_YO �OM_;_q___�_�_�_ �__�_1_�_%ooIo 7omo[o}o�o�_�o	o �o�o�o!E3i �o��Y{U�� ���A��h��1� �������������� [�@��	�s�a����� �������3��W�� K�9�o�]��������� ��/�ɯ#��G�5� k�Y���ѯ������ {�����C�1�gϩ� ��ͿW��ϯ������� �	�?߁�fߥ�/ߙ� �߽߫��������Y� >�}��q�_���� ������������� 7�m�[���������� �����!3i W������}�� �/e�� �U����/� /m�d/�=/�/�/ �/�/�/�/?E/*?i/ �/]?�/m?�?�?�?�? �??OA?�?5O#OYO GOiO�O}O�O�?�OO �O_�O1__U_C_e_ �_�O�_�O{_�_�_	o �_-ooQo�_xo�oAo co=o�o�o�o�o) koP�o�q�� ����C(�g� [�I��m�������ُ � �?�ɏ3�!�W�E� {�i�����؟��� ���/��S�A�w��� ��ݟg�ѯc����� +��O���v���?��� ��Ϳ��ݿ��'�i� Nύ�ρ�oϥϓ��� ������A�&�e���Y� G�}�kߡߏ������ �ߵ��߱��U�C�y��g���������$�SERV_MAI�L  ���~��OUTPUT����RV 2�؍�  � (����_���SAVE����TOP10 �2�9� d  	��������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/�}/�/�/�/���YP�|���FZN_CF�G ڍ����j��!GRP� 2��'&� ,�B   A=0��D�;� B>0� � B4��RB{21l�HELL�"C܍�$�L�M�7|�?�;%RSR�? �?�?O�?%OOIO4O mOXOjO�O�O�O�O�O��O_!_3^�  �R3_a_s_AR_� ��{_�R�P)�xWIR2��d�\�]|�Rh6HK 1�v; �_o"ooFo oojo|o�o�o�o�o�o �o�oGBTf~b<OMM �v?��g2FTOV_E�NB��A�$��ROW_REG_UI����IMIOFWD�L�pߥ~@5�WAIT�r�Y�8��r�v@�0�TIM�u7��j�VA��A�>�_UNIT�s��v$�LC�pTRY�w�$���MON_�ALIAS ?e�yH�he��%�7� I�[�i�������� m����
��.�ٟR� d�v�����E���Я� �����*�<�N�`�� q�������̿w��� �&�8��\�nπϒ� ��O���������߻� 4�F�X�j�ߎߠ߲� ���߁�����0�B� ��f�x����Y��� ��������>�P�b� t�������������� (:L��p� ���c��  �6HZl~)� �����/ /2/ D/V//z/�/�/�/[/ �/�/�/
??�/@?R? d?v?�?3?�?�?�?�? �?�?O*O<ONO`OO �O�O�O�OeO�O�O_ _&_�OJ_\_n_�_�_ =_�_�_�_�_�_�_"o 4oFoXooio�o�o�o �ooo�o�o0�o Tfx��G�� ����,�>�P�b� ���������Ώy�����(�:���$S�MON_DEFP�RO ����c� �*SYSTEM�*M�RECALL� ?}c� ( �}A���şן���� ��2�D�V�h�z� �����¯ԯ���
� ��.�@�R�d�v���� ����п���ϙ�*� <�N�`�rτ�ϨϺ� ������ߕ�&�8�J� \�n߀�ߤ߶����� ���ߑ�"�4�F�X�j� |��!���������� ���0�B�T�f�x��� ������������� ,>Pbt�� �����(: L^p���� �� /�$/6/H/Z/ l/~//�/�/�/�/�/ �/?�/2?D?V?h?z? �??�?�?�?�?�?
O �?.O@OROdOvO�OO �O�O�O�O�O_�O*_ <_N_`_r_�__�_�_ �_�_�_o�_&o8oJo�\ono�ol+cop�y mc:dio�cfgsv.io� md:=>19�2.168.56�.1:10496��o�o�oi5�bf�rs:order�fil.dat �virt:\temp\�o�ogy�:a-#v*.d7I}�Q���fxy�zrate 61 ��q��f�x���b�8#5xmpbac�k�U����� }-/�cdb�p*��ʏ`ӏd�v�����3x��:\,���>�Y�W��(�����4��a���� T�؟i�{�������;� V��������B�ԯ e�w�����/�A�ҟ� ��������P�a�s� �Ϙ���3�ί����� �(���L�]�o߁ߏ���$SNPX_A�SG 2�������� 7 0��%������  ?���PAR�AM ��^�� �	��P��e����*�����OFT_KB_CFG  �ô՞��OPIN_SIMW  ��%�������RVQS�TP_DSBk��%����SR �>�� � &)�%������TOP_O�N_ERR  �/�W�L�PTN ����A�H�RING_PR�MV� ��VCNT_GP 2��'��x 	������`�� ��$��VD��RP 1���(� ��_q��� ����%7 I[m����� ���/!/3/Z/W/ i/{/�/�/�/�/�/�/ �/ ??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_r_o_�_�_�_�_ �_�_�_�_o8o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c����� ������Ϗ���� )�P�M�_�q������� ��˟ݟ���%�7� I�[�m��������ܯ�ٯ����!�3�=P�RG_COUNT�L���[�_�EN�B��Z�M��N䑿_�UPD 1��T  
H���ۿ� ��(�#�5�G�p�k�}� �ϸϳ����� ���� �H�C�U�gߐߋߝ� ���������� ��-� ?�h�c�u����� ��������@�;�M� _��������������� ��%7`[m ������� 83EW�{� �����/// //X/S/e/w/�/�/�/ �/�/�/�/?0?+?=?�O?x?s?�?Q�_IN�FO 1�ɹ�� �F��?�?�?O�9����aA�>>�O�?�1���>O\�YSDEBSUGi�ʰ�0d���z@SP_PASS�i�B?�KLOG� �ɵ��r�0eH�?  �����1UD1:\x�DiO�A_MPC�M�ɵ:_L_ɱ�Aj_ �ɱVSAV �`�MA�A�B�5 X�SVnKTEM_T�IME 1��G.�� 0�0!�4�U�oQ�T1SVGU�NSİj�'����`ASK_OPT�IONi�ɵ�����?a_DI�@��[eB�C2_GRP 2��ɹ�U�o�0@� � C��clBCC�FG �k�\ 9QO
~`
EO B-Rxc��� ������>�)� b�M���q��������� ˏ��(��L�7�p����4m���n�ϟ� \�����;�&�_�q^ �QdT�������ѯ�� �����)�+�=�s� a���������߿Ϳ� ��9�'�]�Kρ�o� �ϓϥ����Ȭ���� �1�C���g�U�wߝ� �������߳�	���-� �Q�?�a�c�u��� ���������'�M� ;�q�_����������� ����7��Oa ��!���� �!3EiW� {�����/� ///S/A/w/e/�/�/ �/�/�/�/�/??)? +?=?s?a?�?M�?�? �?�?O�?'OO7O]O KO�O�O�OsO�O�O�O �O_�O!_#_5_k_Y_ �_}_�_�_�_�_�_o �_1ooUoCoyogo�o �o�o�o�o�o�?! ?Qc�o�u�� �����)��M� ;�q�_�������ˏ�� �ݏ��7�%�G�m� [��������ٟǟ� ���3�!�W�o��� ����ïA��կ��� �A�S�e�3���w��� ��ѿ������+�� O�=�s�aϗυϧ��� ��������9�'�I� K�]ߓ߁߷�m����� ���#��G�5�W�}� k����������� ��1��A�C�U���y� ������������- Q?uc��� ������/A _q�������/� �$TB�CSG_GRP �2����  �  
? ?�  J/\/ F/�/j/�/�/�/�/�/��/;#"*#�1,d�0?1?!	� HD 6@�Y3>��5O1B�H!x?�9D)��6L�ͣ1>���g6�0C�?�?�?�>p�?MCj���?5GB�B��OO)HY�0|Afff?IC�]O_O)O�2 �It?�N\0�/ XU&_ �O_Q_n_9_K_�_�_��[?��C �!�	�V3.00�R	�rc65�S	*`�T"o�V�4�T�p�Y G`mHo + � ��@�_�o��c#!J2*#�1-��o�hCFG ���;!C!�j�rB"]o~� BPz�Pva�� �������<� '�`�K���o������� ޏɏ��&��J�5� n�Y�k�����ȟ��� ���\	��-�ן`� K�p���������ޯɯ ��&�8��\�G��� k�����!/ۿ�� ���5�#�Y�G�}�k� �Ϗϱ���������� �C�1�S�U�gߝߋ� �߯�����	����?� -�c�Q���Y���� m������)��M�;� q�_������������� ����%I[m 9������� !E3iW�{ �����/�// /?/A/S/�/w/�/�/ �/�/�/�/?+?��C? U?g??�?�?�?�?�? �?�?OO9OKO]OoO -O�O�O�O�O�O�O�O _�O!_G_5_k_Y_�_ }_�_�_�_�_�_o�_ 1ooUoCoyogo�o�o �o�o�o�o�o	+ -?uc���� y?����;�)�_� M���q�������ݏ� ����7�%�[�I�� ������o�ٟǟ��� �3�!�W�E�{�i��� ������ï����� A�/�e�S�u������� ���ѿ�����+� a��yϋϝ�G��ϻ� �����'��K�9�o� �ߓߥ�c��߷����� ��#�5�G���}�k� ������������� �C�1�g�U���y��� ��������	��- Q?a�u��� ����/��� q_������ �/%/7/�/m/[/ �//�/�/�/�/�/? �/?!?3?i?W?�?{? �?�?�?�?�?O�?/O OSOAOwOeO�O�O�O �O�O�O�O__=_+_ M_s_a_�_C�_�_ }_�_�_o9o'o]oKo �ooo�o�o�o�o�o�o �o#Yk}� I������� ��U�C�y�g����� ����я����	�?� -�c�Q�s�u������� �ϟ��)�;��_S� e�w�!�����˯��ۯ ݯ�%��I�[�m���=�����ǿ���վ s �� ��)���$TBJO�P_GRP 2��ݵ� / ?��	A�H���O��� ����p{Xd� ���� � �,�� @�`�	 ߐD ��C?aD���`�x�¹���>���ϼ����<!a���?�����>L��?B�  B��8��C�D)�U�CQ?p�D�S�����>���u߻�ff�f���\<��Y�U��C +Р/�<��S�D5m�Κ��݁�&�)�333<���U�>���/>��C�й�<��b�Cj��u�b�����a�;�9b�B�!�?8Q��pG�Hc���s����Y��*��&�8��;��6��%�>u[%�DG���� ������*��8�&�<Z;u����� ����S�E/=k �w1����� ,�KeO]�d������ ��	V3.00f��rc65e�*� e��/ ' �F�  F�� �F� F�  �G� GX �G'� G;� �GR� Gj` �G�� G�| �G� G�� �G�8 G�� �G�< H� ?H� H��2 �Ez  E�@ _E�� EB F� �FR FZ F�� F� F�P<"G � GpL#�?h GV� G�nH G�� G��� G�( =^b�=+�8�$E�Q�?2�=3?�  ��M?�[:A��*SYS�TEM
!V8.3�0218 �38/�1/2017 �A y�p7M�T�P_THR_TA�BLE   $w $�1ENB��$DI_NO��O$DO�4���1�CFG_T � 0�0MAX_I�O_SCAN�2M;IN�2_TI�2D;ME\��A�0�  � $�COMMENT �$CVAL�	CT�0PT_ID�X��EBL�0NUMQBENDIJfAZI�TID]B $DUMMY13���$PS_OVE�RFLOW�$��F�0FLA�0Y�PE�2�BNC$GLB_TM�7�EF@��1�0ORQCTR�L�1 X $�DEBUG�CRP��@2@  $S�BR_PAM21�_VP T$S�V_ERR_MO�DU4SCL�@RA�CTIO�2�0GL�_VIEW�0� 4 $PA$UYtRZtRWSPtR^�A$CA@A�1��1aQUeU �0N�P3@$GImF3@}$eQ lP8_S�PiQ LpP�V�I<P�PF�RE�VNEARPLAN�A�$F	iDIST�ANCb�1JOG�_RADiQ�0$JOINTSP� 	RE_SMS�ETiQ  �WE<�UACONS2@�0��TONFiQ	�? $MOU1A`��$LOCK_F�OL�A�2BGLV�@CGL�hTEST�_XM@@raEMP�E`,R�b�B`�$cUS;AfPH`2Pt�S�a�bMP_�`z�aQCENEdR~r $KARE�@}M�3TPDRAhP|;t2aVECLE�3�2dIU�aqHE�`TOOLH`�0qs�VI{sRESpIS�32�y64�3ACiHX`�`~qONLE��D29�B�pI�1�  @$RAI�L_BOXEHa�PROBO�d?�~QHOWWAR�0x�r�@�qROLM�B2�A�C �SK�r�@n�0O_F9�!�H�S�qiQ
>n�0RVp�OCiQ>bSLO�GaK��VOUZb�R�eAELEC�TE<P`�$PI=P�fNODE�r�r��qIN�q2^��pCORDED�`�`}��0P9P@  wD �@OBAU`TA�a����C�@��p�P�q0��ADRAܥ0F@TCHup 7 ,�0EN�2�1A�a_�Tl�Z@�BޣRVWVA!A� � ApeR�5P�REV_RT�1�$EDIT��VS�HWR9�S@	UАI�S`yQ$IND�0@1QB蓗q$HEAD�5@ ��p5@溒KEyQ�@CPS�PD�JMP�L��5�0RACE�4U�a�It0S�?CHANNEzp��	WTICK{s�1M�`A�0@�HN�A�D0^�]D�`CG�P8���v�0STYf��q�LO�A�SB���jP� t 
��Gr�%�$���T=PS�!$UNIGa5A�E��0�FPORT��SCQU5ptR���B��TERCJ@*b�T=SG� �PPL6�$�DE��$`Thqb�0OK@>CV�IZ�D4�Q�E�APR�A�Ͳ�1��PU}aݵ_�DObk�XSV`KN�6AXI��7�qgUR_s�E$T�p���*��0FREQ_,hp<�ET=�P�b�OPARA`@.P
@�:[���ATHr�3@a�D�s�s�0 .��p�R_Q�0l8}��@�1TRQIc���$`�@��BRup��VyE@@��NOLD��AAp7a��x@�A��AV_MG����¨/���/�D)�D;�D�M�J_ACC.�C��<�CM��0CYC0M@3@��M@_E������٘@o�TSS}C�@  hPcDS���1�@SP�0*�AT:����@��i�~�BADDRES{s=B��SHIF}b�aK_2��S@��I�@�|��TV�bI�2�]��h>��C�
�j
�RV����0 \��������웱�@��CnӞ�aºꯆ:R����TXSCREE���0�TIN!AWS�P;��T�1>�>�jP TQ�7P�B �6QP��
��
�>��RROR_"a�@����D�QUEG�# ���U��@SXQ��RSM�� �UNEaXg��6��0S_�S���	0��>�Cx�b��o� 26�UE���2GRU�ͰGMTN_FL�Q�#POi�BB�L_�pWg@�0 �����O�Q�L1En���pTO`C��RIGH�BRD<ITd�CKGRg@��TEX,���WIDTH�sݐB�A�AZ{q��I_/@H�� � $LT!_ �|�Y0@RyP�b �s�w�B��GOu��0%D0TW� U� �9R�b�LUM�!Ǝ^�ERV��]PFP�`>��1'@r�G�EUR�cF\��Q)&��LP�Z�Ed��)'�$(�$(�p#)U5!+6!+7!+8"�b�>CȰ`��F�qږaS�@EUS=ReT  <��/@qU�R��RFOChq.�PPRIz�m�@?A�� TRIP�qm��UN�0�4!�P  ��0�5�7��b;�5�� "T� ̱G ��T7���}�O2O	SNAd6RA���;3wq�1#n_�S�^�2�����aU!"A$�?�?+8"��;3OFF�` P�%O��3O@ �1#PD,D$PG�UN#K`S�B_�SUBBPk SR	T�0��&��"avp��sOR�p�ERAU���DT�Ib��VCC���H�' ��C3�6MFB1ĢSP=G?�( (b`�STE�Qʀ9PWT�ѠPE���GXd)� ����JMOVE��{Q6RAN4`?[�3�DV�S6RLIM_X �3qV�3qV\XvQk\:`V1�IP�2VF� �C|`�A����*���IB�P,�S� _��`�p�b���@ (0GB�� "P�@��|pr+x �r �,�tRn@��s 9C@TeDRI�PSfBQV!�wdԐ��D�$?MY_UBY�$\d �;QA�S���h�q��bP_S�ף�bL��BMkQ$j�DEYg�EX� ���B_UM_MU6�X�D<q US��?��;V=Go�PACI�TP �<Uyr�3yrkSyr:�;qREnr�1l��8dyr�@,�BTAREGPP�q8eR{0�@- d��;cBi	:r��R�DSWqp$�Sn�:s˰O�!d�QAv�3���E��Up0m��vHK�.��K�AQ��0���?SsEA����WOR�@�3��uMRCVr/� ��O��M�@C��	ÂC�sÂREF��̆��gRj�
� � Ȋ�ي��=�̆r�_RC��s���� �@����b���:bo0 �Т�;��� �e�OU���r��$\c(`+�u��2��<���̰� -=���f�]K�SUL3a.��C7Po/+p�NT�a��]��ag��g��!g�&�L�c���c��(����!�@T�����1���o@AP_�HUR�ۥSA>SCMP��F�����_&�R�T�������X.���GFS�E2/d �M� � Y0UF_�����J��RO� ����W,rUR�GR�mq�AI���D_V_h[D�@�zY��3�WIN.rH���X-V
A�RqR�P�WEw�w�q|c6v�,q��RvLOiPtc��Ld��3t m+=�PA' =�CACH6����ŵ��,p����K�ۓC�QIo�FR"�T� $֭�'$HO�@�R��`� rc��[�֘p��ڔ��VP�r����_S�Z3p���6����1�2� ��]p�؆P��W�A3�MP��aIM5Gx���AD�q�IMREٔ6�_SIZ�P��!po�6vASYNBUF6vVRTDh�t�F�?OLE_2D�T��t��0C0aUs��Q�P�X�ECCU�xV�EM�p����#�VIsRC��VTP������G�p��t��L�A�s�!��qMco4���;�CKLAS�QC	��ђ�@5  ��A�� @&B�T$8��$`��6 |F@o���Xñ�T�o�?a���"�uI���r/��`B�G� VEJ�`PK�|p1�1֖G�_HO|+��R7 � }F����ESLOW�}w]RO>SACCaE*@-�=�xVR:�0�11�yrAD�/0FrPA��&�D�1��M_Ba� ���_JMP���A8|y�b�$SSC6u ��M��C��@92���S8��N/�PLEX��: T〲C�Q���6�FLD?1DEZ�FIQ rO�q�ty�F��PP2��;O� ϱPV�>��MV_PIZ���G�BP��`а�FIQ�PZ�$���0����GA%p��LOO0Tp�JCB�T*����� ��ړPLCAN�R&�L�F�� �cDV�'M�p���U�$�S�P.q�%�!��%#�㱶C4G�����RKE�1�V�ANC]G�A0p �<�@�?�?J�R;_A�a =�?q?�?T0�9���r> hܰ�	��K9�fA2b�<X@̠OUe�ݒA���
O���SK(�M��VIE�p2= �S0:�|R? <�{@XMԊ`UMMYR����Re��D����X�CU��`b�U�@@ $��@TIT 1$�PR8�UOPT?�VSHIFʀ�A`�a���T�0l����$�_R$�UړQ.qZ�U�s�o�t�Qav�Q5fST�G@cVSCO��vQCNT���3� }w�RlW �RzV�R�W�R�XLo^oTpjjA2��51D>a��0� �pSMEO��B%X�J�@�1u���_���@C4%�Gi�LI� ��^'��XVR�DDY���@T� �ZABCP�E�r�bMӺ�
�1ZIP�EF,%��LV��L���}J�ZMPCF�eMGy�$p?�r?DMY_LN$@A8r8��dH ���g�\�>�MCMİC�ӟCART_Xq�P~�1 $JvsptD��|r�r�w���u����UXW�puU�XEUL�x�q�u �t�u�q�q�y�q�v r�eI Hk�d����Y�`D�� J� 8o�	V�EIGH��H?("��f�9�ĔK �= �C,���`$B&�K���1�_�B��LgRV� F8^���COVC؀qr@fq9��@}�e�
��4��7�D�TRȰ?�9V�1�SPH� ǑCL !�S�i�{�����ST�S  g������0��0�u�<�ѐNa1 ��;�� ����T����������U��������	���a�����������������1��'RDI������ğ ֟����t�O|���@������ίஔ�Sz��� >�����ſ׿� ����1�C�U�g�y� �ϝϯ���������� v�}���8�!�3�E�W� ��'�9�K�]���Ҷ ����
U�5` Y��0�����0��@A�v�^`BF_TT��ի���BI�V>0�2J�_�I��R 1&� 8!����%к� ��C�  ����������� �"�4�F�X�j�|��� ����������1�gBTjx�� ���р����0B QI�Zl J�������� �/"/4/F/X/FҒ� t/�/b*���/�/��b�v�@`�v�MI_�CHANU� `� �#3�dV�`�u�&0E}T>�AD ?��y0�m��/�/�?Ȥ?�d0RLPs�!�&�!�4�?�<SN�MASKn8��1/255.4E0�33O�EOWO�OOLOF�S^Q �`�$X9OR�QCTRL D&�V�m��O��T�O �O
__._@_R_d_v_ �_�_�_�_�_�_�_o�o(l�OKo:ooo��P�E�pTAIL8�JP�GL_CONFI�G 	�ᄀ�/cell/$�CID$/grp1so�o�o1�#��?\n���� E����"�4�� X�j�|�������A�S� �����0�B�яf� x���������O���� ��,�>�͟ߟt��� ������ίB�}c�� �(�:�L�^���`o��e��b���Ϳ߿�� �\�9�K�]�oρϓ� "Ϸ����������#� ��G�Y�k�}ߏߡ�0� �����������C� U�g�y����>��� ����	��-���Q�c� u�������:������� );��_q� ���H�� %7�[m�����]`�Us�er View ��i}}1234567890�
//�./@/R/Z$� �cz/���2�W�/�/�/@�/??u/�/�3�/ d?v?�?�?�?�??�?�.4S?O*O<ONO`OrO�?�O�.5O�O�O��O__&_�OG_�.6 �O�_�_�_�_�_�_9_�_�.7o_4oFoXojo |o�o�_�o�.8#o�o �o0B�ocir� lCamera��o�� ����NE�,� >�P��j�|�������ď�I  �v�)�� &�8�J�\�n������ ���ڟ����"�4�[��vR9˟������ ��ȯگ�����"�m� F�X�j�|�����G�Y� I7�����"�4�F� �j�|ώ�ٿ������ ����߳�Y�����Z� l�~ߐߢߴ�[����� ��G� �2�D�V�h�z� !߃unY��������� ����B�T�f���� ������������Y�"i {�0BTfx�1� ����, >P��Y��i��� �����/,/>/ �b/t/�/�/�/�/cu9H/�/?!?3?E? W?�h?�?�?F/�?�?@�?�?OO/O�j	�u0�?jO|O�O�O�O�O k?�O�O_�?0_B_T_ f_x_�_1OCO�p�{._ �_�_oo+o=o�Oao so�o�_�o�o�o�o�o �_�u���oOas ���Po���< �'�9�K�]�o�PE c����͏ߏ��� �9�K�]��������� ��ɟ۟����ϻr�'� 9�K�]�o���(����� ɯ�����#�5�G� �;�ޯ������ɿ ۿ���#�5π�Y� k�}Ϗϡϳ�Z����� J����#�5�G�Y� � }ߏߡ�����������x����  �� N�`�r��������������    $�,�J�\�n������� ����������"4 FXj|���� ���0BT fx������ �//,/>/P/b/t/܆/�  
��( � �B�( 	 �/�/�/�/�/?? 8?&?H?J?\?�?�?�?�?�?�*4� � n�O1OCO��gOyO�O �O�O�O��O�O�O_ VO3_E_W_i_{_�_�O �_�_�__�_oo/o AoSo�_wo�o�o�_�o �o�o�o`oroO as�o����� �8�'�9��]�o� ���������ۏ��� F�#�5�G�Y�k�}�ď ֏��şן����� 1�C�U���y������ ��ӯ���	��b�?� Q�c�����������Ͽ �(�:��)�;ς�_� qσϕϧϹ� ����� �H�%�7�I�[�m�� �ϣߵ��������� !�3�E�ߞ�{��� ������������d� A�S�e���������� ����*�+r�O�as������0@� �������� ��)frh�:\tpgl\r�obots\r2�000ic6_165f.xml� `r�������/����/3/E/ W/i/{/�/�/�/�/�/ �/�//
?/?A?S?e? w?�?�?�?�?�?�?�? ?O+O=OOOaOsO�O �O�O�O�O�O�OO_ '_9_K_]_o_�_�_�_ �_�_�_�__�_#o5o GoYoko}o�o�o�o�o �o�o o�o1CU gy������ �o��-�?�Q�c�u� ��������Ϗ���K � 8?8�?��2� �.�P�R�d������� ���П���(�R��<�^���r�����ܫ��$TPGL_OUTPUT ���� � ���%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ�������ˠ2345678901�� ������0�8����� _�q߃ߕߧ߹�Q߽�@����%�7���}A� i�{����I�[��� ����/�A���O�w� ��������W����� +=����s�� ���e�' 9K�Y���� �as�/#/5/G/ Y/�g/�/�/�/�/�/ o/�/??1?C?U?�/ �/�?�?�?�?�?�?}? �?O-O?OQOcO�?qO��O�O�O�O�OyO֡} �_)_;_M___q_�]�@��_�_� ( 	 ���_�_o �_5o#oYoGoioko}o �o�o�o�o�o�o /UCyg��� �����	�?�����-�G�u���c��� ����ߏ���`��,� ΏP�b�@�������� Οp�ޟ����:�L� ��p���$�������ܯ �X���$�Ư�Z�l� J������ƿؿz��� ��2�DϮ�0�zό� .ϰ��Ϡ�����b�� .���R�d�B�tߚ�� ����߄�����<� N��r��&���� ����Z�l�&�8���\� n�L����������|� ���� FX��| �0�����d 0� fxV� ����//� >/P/�</�/�/:/�/��/�/�/?
2�$T�POFF_LIM� [��@W�y��A2N_SV#0�  �T5:P_�MON S�)74�@�@2�U1�STRTCHK �S�56_=2VTCOMPATJ8��196VWVAR �j=�8N4 ��? O�@}2�1_DEFPRO/G %�:%&OmO�;4_DISPLA�Y*0�>?BINST�_MSK  �L� {JINUSE9R�?�DLCK�L�K�QUICKMEN��O�DSCREP�S��2tps�c�D�A1P6Y52GP_�KYST�:59RACE_CFG �F�r1�4.0	D
�?��XHNL 2E�93��Q�; $B �_�_o o2oDoVoho�zj�UITEM 2��[ �%$1�23456789y0�o�e  =<�ox�o�os  !{!@�oZC�o{ �o���9K� o/��?�e���� ��#���G���+� ��O���ŏ׏Q����� ͟ߟC��g�y���� ]������������-� ��Q��u�5�G���]� ϯ!����ſ)�տ�� �q�ϕ�����3�ݿ �ϯ���%���I�[�m� ��	ߣ�c�u��ρ��� ���3���W��)�� ?���ߌ��ߧ��� ��c�S�e�w���� ��k��������+�=� O���s�EW��c ������9� o��n��� ��#�G�"/} =/�M/s/�/��// /1/�/U/?'?9?�/ ]?�/�/�/i?�??�? �?Q?�?u?�?PO�?kO �?�O�OO�O)O;O_ʐTS�R�_UJ�g  �bUJ �Q`_UI
 m_�_z_��_8ZUD1:\��\��QR_GR�P 1�k� 	 @`@o!k�oAo/oeoSo�own� �`�o�j�a�_�o�o�e?�  '9{# YG}k���� �����C�1�g�U�w���	�E��Ï~SSCB 2%[ �!�3�E��W�i�{�����\V_�CONFIG �%]�Q]_�_���O�UTPUT <%Y�����S� e�w���������ѯ� ����+�_A@�S�e� w���������ѿ��� ��+�<�O�a�sυ� �ϩϻ��������� '�8�K�]�o߁ߓߥ� �����������#�5� F�Y�k�}������ ��������1�B�U� g�y������������� ��	->�Qcu ������� );L_q�� �����//%/ 7/H[/m//�/�/�/ �/�/�/�/?!?3?D/ W?i?{?�?�?�?�?�? �?�?OO/OAOݟ� >�O�O�O�O�O�O�O �O_!_3_E_W_J?{_ �_�_�_�_�_�_�_o o/oAoSod_wo�o�o �o�o�o�o�o+ =Oaro���� �����'�9�K� ]�n��������ɏۏ ����#�5�G�Y�j� }�������şן��� ��1�C�U�g�x��� ������ӯ���	�� -�?�Q�c�t������� ��Ͽ����)�;� M�_�p��ϕϧϹ��� ������%�7�I�[� m�~ϑߣߵ������� ���!�3�E�W�i�LH������� s���hO������1� C�U�g�y��������� t�����	-?Q cu������� �);M_q �������/ /%/7/I/[/m//�/ �/�/�/��/�/?!? 3?E?W?i?{?�?�?�? �?�?�/�?OO/OAO SOeOwO�O�O�O�O�O �?�O__+_=_O_a_ s_�_�_�_�_�_�O�_ oo'o9oKo]ooo�o �o�o�o�o�o�_�o #5GYk}�� ����o���1� C�U�g�y����������ӏ���$TX_S�CREEN 1������}��&�8�J�\�n���������ҟ� ��������P�b�t� ������!�ίE��� �(�:�L�ïp�篔� ����ʿܿ�e�w�$� 6�H�Z�l�~������ ��������� ߗ�D� ��h�zߌߞ߰���9� K���
��.�@�R��� v��ߚ����������k���$UALR�M_MSG ?��� ��zJ� \��������������� ����/"SFw+��SEV  �E���)�ECFG ���  }�u@�  A��   B��t
 x�s�0B Tfx�����~�GRP 2�w 0�v	 ��/+�I_BBL_NOTE �
�T��l��r��q� +"DE�FPRO5�%9� (%k�/�p�/�/ �/�/�/?�/%??6?�[?F??j?�?!,INUSER  o-�/�?I_MENH�IST 18�� � (�  ���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1�?`OrO�O�O�s� (O:M936MO �O�O__�B/_A_S_ e_w_�_�_*_�_�_�_ �_oo�_=oOoaoso �o�o&o�o�o�o�o '�oK]o�� �4�����#� �<V""A�_�q����� �����ݏ���%� 7�Ə[�m�������� D�V�����!�3�E� ԟi�{�������ïR� �����/�A�Я� w���������ѿ`��� ��+�=�O�:�L��� �ϩϻ�������� '�9�K�]��ρߓߥ� ��������|��#�5� G�Y�k��ߏ����� ����x���1�C�U� g�y������������ ����-?Qcu `�rϫ���� );M_q� �����//� 7/I/[/m//�/ /�/ �/�/�/�/?�/3?E? W?i?{?�?�?.?�?�? �?�?OO�?AOSOeO wO�O�O���O�O�O __+_.OO_a_s_�_ �_�_8_J_�_�_oo 'o9o�_]ooo�o�o�o �oFo�o�o�o#5 �o�ok}���� T����1�C���g�y����������O���$UI_PAN�EDATA 1������  	�}ӏ��,�>�P�b�t� ) v���V��şן��� ����C�*�g�y�`� �����������ޯ���?�Q�8�u�R�� �A������Ŀֿ ����_�0ϣ�B�f� xϊϜϮ���'����� ����>�%�b�I߆� ��߼ߣ����������7���T�Y�k�}� �������J���� �1�C�U���y���r� ����������	��- QcJ�n�� 0�B��);M �q������ �/h%//I/0/m/ /f/�/�/�/�/�/�/ �/!?3??W?���? �?�?�?�?�?:?OO �AOSOeOwO�O�OO �O�O�O�O�O_ _=_ O_6_s_Z_�_�_�_�_ �_�_d?v?4O9oKo]o oo�o�o�_�o*O�o�o �o#5�oYkR �v������ �1�C�*�g�N����� o"oӏ���	��-� ��Q��ou��������� ϟ�H���)��M� _�F���j�������ݯ į����7�����m� �������ǿ���� p�!�3�E�W�i�{�� �φ����ϼ������ /��S�:�w߉�p߭�0����D�V�}���� -�?�Q�c�u�)	�� ŉ���������� � ��D�+�h�O�a����� ����������@�R9v	�`�Z��$�UI_POSTY�PE  `�� 	 ����QUICKM_EN  ����� RESTOR�E 1 `�  �iB�S`N�m~ ������/%/ 7/I/[/�/�/�/�/ �/r�/�/�/j/3?E? W?i?{??�?�?�?�? �?�?�?O/OAOSOeO ?rO�O�OO�O�O�O __�O=_O_a_s_�_ (_�_�_�_�_�_�O�_ o"o�_Fooo�o�o�o �oZo�o�o�o#�o GYk}�:o�� �2���1�C�� g�y���������d�����	��-��SCR�E� ?��u1scHu2�h�3h�4h�5h�6�h�7h�8h��US#ERJ�O�a�TI�j�Sksr�є4є5є�6є7є8ё� N�DO_CFG �!����Ѩ PDA�TE ���None _� ���_INFO 1e"`�]�0%3� x�	�f�����˯ݯ�� ����7��[�m�P��������ǿ�J�OFFSET %�ԿσA֏�*�<� N�{�rτϱϨϺ�� �����A�8�J�w�@n߀ߒ�����
�����UFRAME�  ʄ�G�R�TOL_ABRT8&��>�ENBG�8�?GRP 1&<Cz  A��� ���������������:�� Ug��V�?MSK  j�]�JX�N#���]�%�߼���VCCM�Y'���RG��*�	Q��ʄƉD � BH)�p<2Ce�)��PN?�` 6��MR��20��p���"�р	 ���~XC56 *�d�����N�5рm�A@<C�' ���ʈ�);h�c���Rр|�Ђ? B����6 �t/T1/ /U/@/ y/d/�/�/�/�/*/�/ 	?�/???�c?u?��TCC��1��f�9��рр��GF�S�22w ����2345678901�?�2ʈ"�6� �?!Oс>,12�QO_G�B@R 8N:�o=L���� �������OOA�O �O@O_dOvO�O�O�O �_�O�O�___�_<_ N_`_r_Soeo�_Ro�o �_�_oo&o8o��4SELECF�j��$�VIRTS7YNC� ��6��BqSIONTMOiU-tр��cu���3U��U��(�� FRk:\es\+�A\�o� �� MC�vLOG�   oUD1�vEX��с' B@ ����q�o6��q�:�^�σ � � =	 1- �n6  -���ʆ�xf,p�#�0=���ʹ���r>�xTRAIN��2(�1.��
. d��s:q4w (,1�� 0��)�;�M�_�q��� ������˟ݟ����I��crSTAT 5��@%������E:$��ۯ�_GE���6w�`. ��
��. 2�HOM�IN��7U��U� �r�a�a�a�CG�um�JMP�ERR 28w
  ʯE:��suTs �����߿���'π9�O�]ώρϓ�_v_��pRE��9t���L�EX��:wA1-�e�VMPHASOE  RuCCb���OFFLpc�<vPU2�t;4�04��8�
��b@�� �bb>?s33��Á�1��L��ҕԈ�|��
t�>x��Â�xf�o�.���/?P�X�  $�2�x����0� � ��6�+���l��\� j�|���������� � D�V���ZTf� ���������.  �,BPb��� ����//(/ :/�y/�b/��/� /L/? ??<?n/c? �/�/�?�?�/�?6?�? �?�?OX?j?\O�?�O JO�?fO�O�O�O�O0O %_TO_xOm_�O�O�O �_�_�_�__o>_P_ EoWo�_xo�_�o�o�o��o��TD_FIL�TEt�?�� ��Wp��]o$6H Zl~����� ���)�;�M�_��q������SHIF�TMENU 1@x�<��%���� я��0���f�=�O� ��s�����䟻�͟����P�'�	LIVE/SNAPD�vsfliv��b���ION� G�U���menu����:�����±�6��A���	����Lb�K��5M����m`�@�����A�pB8
������Ӝѝ���9���m`� ;ӥ��/�ME��uY��ZM���MO��B����z��WAITD_INEND�3����OKN�.�OU�T#��Sa�4�TI]M�����G� ��@���`ϱ�ϱʞ��2�RELEASE�����TM���=��_ACTx������2�_DATA C�ի�%i��ߪ����RDIS�b�_�$XVR2�D���$ZABC_G_RP 1E8�n`�,@h2��ǽZIP1�FD� cCo�������x�MPCF_G 1G8�n`0<o ����=�H8����t� �	�w�  8�R�����e�����?� k������5��
\���  � a �����7������I��z��YL�IND�aJ�� ��f ,(  *s�K�p���� �//+.m N/�r/Y/k/�/��/ �/�/3/?�/�/J?1?�n?U?�/�?�?v�C�29K8��� ��O `o�7O~[Ol�?�O�g��AA�ASPHERE 2LS�?�OX?�O__>_ �?�Ot_�_?�_I_/_ �_�_o�_]_:oLo�_ �_�o�_�o�o�o�o#o� $7�ZZ� �k�