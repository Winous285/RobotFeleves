��  gb�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A(  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�   � �ALRM_R�ECOV�  �� ALM"ENB���&ON&! M�DG/ 0 $DEBUG1A�I"dR$3AO� T�YPE �9!_I�F� P $�ENABL@$QL� P d�#U�%�Kx!MA�$L4I"�
� OG�f �d PPINFwOEQ/ ��L A �!�%/� H� �&�)EQUIP 2� �NAMr �'2_�OVR�$VE�RSI3 ��!CO�UPLED� �$!PP_� CES0s!_81F3K2> ��! � $�SOFT�T_I�Dk2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5Xk2S�CREEN_(4n_2SIGE0_?|q;�0PK_FI� �	$THKY�GPANE�4 ~� DUMMY1d�DDd!OE4LA!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTc@�D5�F6�F7�F8�F9�G0�G�GJA �E�GbA�E�G1�G T�F�G1�G2�B �SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HO30IO�0� }%�SMACRO�ROREPR�X� D+��0��R{�T UT�OBACKU��0 �)DE7VIC�CTI*0�A� �0�#�`B�S�$INTERVA�LO#ISP_UN9I�O`_DO>f7�uiFR_F�0AI�N�1���1c�C�_WAkda�jOF�F_O0N�DEL��hL� ?aA�a1bc?9a�`C?��P��1E��#sATB��d��MO� �cE' D [M�c���^qREV�BI�Lrw!XI� QrR�  � OD��P�q$NO�^PM�Wp�t�r/ "�w� �u�q�r�0�D`S p �E RD_E�pCq�$FSSBn&$CHKBD_SE^e�AG G�"$SLOT_��2=�� 	V�d�%��3 a�_EDIm  O � �"��PyS�`(4%$EP�1��1$OP�0�2��a�p_OK�UST1P_C� ��d���U �PLACI4!��Q�4�( raCOM9M� ,0$D�����0�`��EOWBn�IG�ALLOW� �(K�"(2�0VA�Ra��@�2a�B�L�0OUy� ,�Kvay��PS�`�0M�_O]����C�F�t X� GR�P0��M=qNFL�I�ܓ�0UIRE��$g"� SWIT{CHړAX_N�P]Ss"CF_�G�� �� WARN�M�`#!�!�qPLI��I�NST� CO�R-0bFLTR^C�TRAT�PTE�>� $ACC1a��N ��r$ORIأo"��RT�P_S�Fg CHG�0I���rTא�1�I
��T�XP��� x i#�Q�.�HDRBJ; C�,�2'�3'�4'�5�'�6'�7'�8'�9�s!�qCO`T <�F П����#92��L�LECy�"MULTI�b�"N��1�!쇱�0T_}R ; 4F STY�"�R`�=l�)2`�����`T |� �&$�c�Z`�pb��P�M�O�0�TTOӰ�Ew�EXT����ÁB���"2� ��[0]�}R���8b�}� D"}� ���Q���Q�kc1Ă��^ȇ1��ÂM8���P�� ŋ� L�  ���P���`A��$JOB�n�/�i�G�TRIG�  d�p�߻���@³�7�����9��s_M�b! t�p�F� CNG AiBA� ����M���!��@�p� �q��0��P[`X��i�*�"6����0tB񉠎"J��_)Rz�gC�J��$�*?�Jk�D�%C_�;�P�����0h ��R�t#� �������G���0NHAN�C̳$LGa��B@^a��� �D��A�`��gzRɡ�!���p�DB�R�A�AZ�0KE�LT�Ė��PFCT�&��F�0�P��S	M��cI��1�%  ��% ��R��a����B� S��&���M 0�0{o e#HK~�A^S�����Ԡ۠�t�$�"6SW�CSXC)�?!%��p)3���T�$@��PA�NN&�AIMG_�HEIGHCr�W3IDI AVT�0��}H F_ASPװ��`EXP�1��_�CUST�U��)&��|E\�%�C1�NV _�`�a��' 1\%1y�`OR�c,"��0gsk��PO��LBSYI�G��aR%�`���Pspm��0k�DBP_XWORK��(��$SKP_�`G�D�B<qTRp ) ���P���� �0f�DJ!d/�_CN�0�R�#� �'PL�S�Q��d�s�DKA7WA w'�^A�@NFZpfB�DBU��*�"!P	RS�7�
ЖQ����g+ [pr�$1�$ZϢ�Li9,�v?�3ʠ��-�?�4Cr��.�?�4ENEy���� /�?�3J0R�E`��20H��C�uR+$L,C,$pi3
�? =KINE@�fK!_D�I�RO�` ����ȳqvC��h ��FPAÃ3uR�PRYN�B�MR��U!�vu�CR[@EWM ^�SIGN��A�� .q�E�Q-$P���.$Pp 2�	/ P7�PT2�PDu`L���VDBAR@�GO_AW���Jpp � �DCS�p~Z�CY_ 1����@1<�Q?fIG2
�Z2>fN>�����
��qS&c}P2 P M$��RB?�e�P=hPwg�QBYl�`gyT+1�THNDG�23��KS�SE|�Q���SBL�Y�cc�T�G1sQL�4 H�pZ ���VTOFB�l�FEfA�ǿb�T4qSW5�bDOC���MCS�f�`Z$r��b H� W0��TހeSLAV�16�rINP��f��Ly|qQP�7� $,�S���=��v���uFI��r줭s�c�!��!W1ԭrN�TV'��rV	��uSKIvTE�@W����:�J_� _<�00�SAFE�A��_SV��EXCL�U��B �PDJ L�1�k�Y�d�ƻrI�_V� !PPLY� 0b���DE~w��_�ML2�B $VR�FY_�#��Mk�IOU��憻 0���:�O�P��LS�@jb;�#3572��Sr�� Px%X�{P�hs� ��g 8 @� TA� �qঠ �"�`SGN��96����@�A �����iPt!��s"��~UN�0jdՔ�U���B �@� ���Ȼ ���G1l�OG]I�2: @�`Fؒ���OT�@@�:41�(�774C2�M`N�I�2;�R������A܂q��DAY1#LO�AD�T/4~�;30� ��EF�XI�b< @%1O㠈3� �_RTRQ��= �D�`@��Q@  ��EjP"�㥎�<��B�� 	�@��AMP��]>�a���0��a�8Sq�DU�@q�]��"CAB��?A�f�0NSs���IDI�CWRK�^�� V�W�V_]���> ��DI��q�@� �/.�L_SE2�T ���/�Z`��0��#�E_��u�v�j��SWJ�j� 𲰂�d	���=c�OH�fz�PPJ�v�IR!��B� ��w�d��B"����BASh���  X ���V����?C���Q��RQDW��MS���AX}�8�u�LIFE� �7�A1C�NJ���S��H����Cs�>��C�`QN"�U��OV�� _�HE����SUIP�hbC�� _�Ԅ����_����[Q��Z��W���ו�Tbƌ�XZ$ `1��Y2�F�CM@T��t@�N��p�2r��9A `��P.�HE��SI�Zy֥�u��BN�pU7FFI���p� ��Q/40�<26C3��M�SW9B 8�K�EYIMAG�CTM@A��A�Jr|#>��OCVIET���'C C�V L�t���s?� 	G1� :�D�"pST�!x�0�� 0��Ѡ��|0���EMAIL����@����c`_FAU�L��EH�CCO�U�p}$T@��FO< $���eS]�v��ITvBUF�砤q���T  ���BdC�t����#��SAVb$)�e�A� }���Pi�e@�U�b`_ H���	OT{BH�lcPր(0�
{��AX1#�� �@��_GJ�f1YN)_�� Gj�D�U/0�e��M����T
8�F��ِ�A!�H�(@u���C	_r@�@K�D�����=pR���uDS�P �uPC�IM@b��J���U�0�ЁEƀ��IP�su2��D���TH0�c���TuA�HSD=I�ABSC�ts��0Vzp*} �$�#��NVW�G�#�$0$� FJ�/d�j��ASC��U�M�ER��uFBCM�P��tETH�!AI6��FU��DU �a�@;⠂CD�O � ����R_NOAU]Tg` J��P�p2��n4ĥPSm5Cʄ�}5CI�.��`k3� =KH *}1Lp��Q��& �I���4#Q�6s��6@ѡ�60��6���67�9�8�99�:J��8�:1�J1J1J1+J1�8J1EJ1RJ1_J2RmJ2�;J2J2JU2+J28J2EJ2RJU2_J3mJ3�:3KBJ3J/�G8J3EJ�3RJ3_J4mB2qESXT�>aLC`�� F�fF�5Q9g�5���FDR�MT��VC��C�wa}"CҗREM,�FAj�O�VM��eA�iTR�OV�iDTm �jMX�lIN�i���j�'IND�`!�
xp /$DG���`�opS�9�D��`RI�V)0Qbj�GEAR��IO0�K�bu�N j�x�.؎��p�qj�Z_MCM>�C���F��UR)2N y,{1��? ���
 ?�pI�?2�qE���q�d`U �0lbO����P�� �RIT5ca%ET�UP2_ P Ѡ#TD= ��C�����qP�J�,�BAC;Q T��$9 O�-)��OG��%E��3e&0IFI��e0��0����PT���F�MR2ieR ivbY�vbLIq ��{g����f���J�b_mAN~F�_F��I4+�M;v`r}DG�CLF��DGDY&��LD�q>t5[�5�S�كk�S��M�� T�FS� l�T� P�)���
�/�$EX_)�@�)�1P�� ��*�3b�5b�s�G�!ieU � p�&2SWKO��DE�BUG�S��0�GRtY�zU�#BKU� �O1�@ O�P�O8��Π0��ΠM�S]�OO��SMz]�Eq��p�Q`_E V �$�X��p�TERM�2�W;����ORI�Ā6�X;�_`�SM�_��$7�Y;�]���TAy�Z;�/�U}PB�[� -���QbV$G���W$�SEGźאELT}O��$USE0NFI����p����`���X$UFR�����q0豈�D5h�OT1Ǵ TA_ �C�wNSTd�PATT!<��Y�PTHJ!B0�En�K0�ART�� ��������REyL��&SHFTF"��_���_SH��M��!B0x� ��n���Z����OVR
#&SSHI����U�2 ��AYLO$ 5I�1�_�d���d�ERV�0*�} ��b?�d���Q����A��RC<
���ASYMh��F�WJ�apE�����f�2�U��d�5����D5��P#Gи!�	�ORd�M��G	R!���\��΢�^������k�] �tE���TOC�1졳q��OP��N Pz�3&1���aO�a�> RE��R�#&OX0��`�e��R]���������e$PW�RSpIM��[�R_���VISy�r����UD�-���� �^>�$H����_�ADDR9fH$�G a�z�s�i1R� .=_ H8�S� ��S��C��C��CS1E�abaHSO0���` $���_D�`���PR��r�HTT� U�TH�a ({0O�BJE1u���$�9fLEP�-=b� � *g!AB%_qT��Sk�#�DBGLV5#KR�L"�HIT�BG�0LO���TE�M4$��b������S�S�p�4JQUER�Y_FLA��f W(YA���c��� 3PU�"B�IO0���4G��H��HB _�IOLN~�d/0�i�C��$SLz�� PUT_�$���Pwp�rwSLA�� e/2�����ӡ��؁I�O F_AS�f��$L��U���#��04�#����,�H�YOgN!'#�UOP�g ` l!9f�b >$�`E&�!��P�����'�!E&�"�&�P_�MEMBk0T 7h X IPz�v��"_#0v����0��pOc6�1w�DSP��' $FOCUSB}Gv�FS�UJhf�i � 60S��JsOG�W2DIS��J7��O��$J8�97��I6!�2�77_LABQ����0��8�1APHI�p�Q�3�7D+�J7JxRA4`P�_KEYp� �KILM�ON�j&`$X�R =0cWATC�H_ �DӘ�U1EL�� �y`B�k �GpG�VP�-ffBCTaR��fB5baLG|�l ��+h�"��LG_SIZ{Y��E�
��F
 �FFD�HI �H�H��F�HM��F�@ ���C5V
�5V
 5V�@5VM�5W�`S)@S�����@Nv1��mx �� ��R��4a�PÀU��Qk�L�S�RDAU�UEA I���R��PGH���AOG�BOO~�n� C-"2�ITGcd���)&REC-jSCRYN)&DI(#S��RG����cl�!#���b�!Sa"Wpkd!�T!#JGM�g�MNCH"FNt�2�fK�gPRG�i�UF�h	��hFWDv�hHL/ySTP�j�V�hĀ�h`�hRS"gyH!�{&C�Es ��!#���g�yUt@�g�¬f|@6#�bG�i�4�PO�JzZeEsMجw82�iEX'TU%I�eIP�cw��c ���c���`�a����s���Jg��KaNO{�A�NA"貇�VAI̵0zCL����DCS_HI��������1O����SI)��9S'��hIGN�@���C�aT����DE�V�wLL�єQ6@B�U𠔠oa@�T6��$�GEM'9FnD���ҡ��pa@�ЅC�!��OS�1��2��3��d_����q �T0v-�p絡.e�IDX����-fL�b�ST�m R�PY0���� _p$E��C����  ����*3���r L*</��Q(6����6�EN 6��Jd?_ s Y��P�$ dKaD� �MCޜRt �T0CL�DPm ��TRQL�I`��e0x�f�FL >1��_����DUA���LD������ORGe0�r���WX������Y���V�O�u �C 	���uu���Si��Tx��00�ްS�>[�RCLMCi���`�{�m[�*�MI���O�v d�Q6�RQz�00�DSTB���Y� ��{a��AX��@�� �EXCE�S�����M��w�T��¹�+���x(��_A�ʊ l�����V�K|�y \�*�2��$MBL�IE��REQUI�R����O��DE�BUES�ML
�M{�zW�.!��B4��i�Y�MN,03�¨�{�R�RkHV�DC�E��TIN3 `!�TR#SMw0p�S�N����p�s<�ՐC�PST� w |h�LOC9��RI� 9�EX��A���:�����ODAQo%}��$@�Q΂MF�A�_���pp�C��P��SUP��*�FX��IGG�"~ �0��MQ@���v�5@� %�����m ��m ����6#D'ATA����E� 1�)�MQ" N�� tV�MDIF)?�!��H���1!x� �Q"ANSW�a�!ܑS�!D�)�����H3Q�$� ?�CU�@V_ >0��&�LO�P$�=ұ���L2������RR2I5��  ��QAX� ?d$CALI��NU�G�2gRIN�p<$RSWq0��K�ABC�?D_J2SE�����_J3v
p1#SP�@6 ��Pp��3��\����J����P�O��IM<��[�CSKP��$H�P�$J�Q[�Q,�6%%6%,'��_AZW��h!EL�����OCMP����1X0cRT�Q�#�1�c@��Y�1��(�0�*Z�$SMG�p�����ERJ*�I-N� ACߒ��5P�b��1�_B�5�42d���14X҆>9DI~!��DH �30���$Vo�Y�$�a$� ��A��<�.A��ňH �$BELy |lH�ACCEL?���8���0IRC_)R��А�ATw�c�O$PS �k�LM�yP D��0G�Q�FPATH�9WG�3"WG3&B��#�_�2��@�AV���C;@�0_{MG|a$DD�A<@[b$FW(���`�3�E�3�2�HDE�K�PPABN.GROTSPEE�B��_8x�,!��DEFg��1~M�$USE_J��Pz�C ���YP��0V� �YN��A�{`uV�8uQMOUf�ANG�2�@OLGC�TINC~���B�D����W���ENCS�����A�2��@INk�I&Be��Z�, �VE�P'b23_�UI!<�9cLOWL�3��pc x��UYfD��p��Y�� ��Uy�C�$0 fMOS`���M�O����V�PERC�H  vcOV�$  �g9��c��\bYĄ��' �"_Ue@0��A&BuLcT����!ec�\j�WvrfTRK�%h�AY�shчq&B�u�s����&l��Rx�MOM |���h�ﰞ ���Ca�sYC���0DU���BS_BCKLSH_C&B��P�f�`�}S�7��RB��Q.%CLAL��b?��pX�Nt�CHKx�H�S�P'RTY����e������_~��d_UM�l�ĉCу�ASCL�ބ PLMT�_L �#��H�E��� ���E�H�-��Q�#p_��hPC�a�hH���ЯEǅCw��X�T�0�GCN_(N��þ���SF�1�iV _RG�e�!��&B���7CATΎSH~�( �D�V��f�'A�	�� �@PA΄�R_Pͅ�s_y�뀎v�`x��s����JG5�6Ф��G`OG���rTORQUQP��c�y�@��0�b�q�@�_W�u�t��!�14��33��33�I*;�II�I�3F�&�������@VC�00���©�1��2�ÿ����JRK����綒 ?DBL_SM�QOMm�_DL�1O�GRV:�3ĝ33ģ3��H_��Z@a�CO1Sn˛ n�LN���� ���ĝ0��� ��e��ʈ�̃��Z���f�M1Y���z�TH��.��THET0beNK�23�3Xҗ3��CB�]�CB�3C��AS����e��ѝ3��]�SqB�3��h�GTS@! QC���'y��'����$DU��;w	�@�Q�����qQ��N��$NE$T�I��H���)I7${0L�AP��y��`�k�k�LPHn�W�1eW�S����� ����W���������{0EV��V��0��V��UV��V��V��V��V�V�H����P��7�����H��H��UH��H�H�O��O��OF	��O��O���O��O��O��O
�O��FW�}��	������SPBALAgNCE�{�LE��H_P�SP1��1���1��PFULC�5\D\��:1���!UTO_��ĥTg1T2��22N�� �2, ����q^<�-B#�qTHpO~ �1$��INSEG�2{aR�EV�{`aDIF�quC91�('o21��dpOB!d�=��w2���7P���LCHW3ARR�2AB���u?$MECH���X�Q�!��AX�qPB�p�&r�~2�� 
�"���1eROB�`C�R r�%��-S0MS�K_�4� P �_OPR�1�2(47Qst1�,`*R(0)c�B�(0|!IN!�MTCOM_C��>�0�  �@0 ~�A$NOREc�2�l ~2� 4��GR��%FLA�!$XYZ_D�A��LP;@DEBUb�2 �0lR�0� (�$mQCODS� ��2�r� �p$BUFINDX*P�0;@MOR3� H%0�p�0��:@��p�QB�"�1ح�NF�TA9Q�#C�rG.B� � $SIMUL����0�As�AsOBJ�E3�FADJUS<�H�@AY_I��xD�GOUTΠ�4�pn�P_FI�Q=8AT#�Y,`W�1P +��PQ+ 9�uDjPF�RI �PUT0�RO��
`E+�Sp�OPsWO��0�,@�SYSBUi� @$�SOP�QBy��ZU<�[+ PRUNn2�UPA;0D�V�"�Q�`a_�@F��PP!AB�!�H��@IMAGS�4%0?�P!IMQAd�IN$��RcRGO�VRDEQ�R�@�QP0�Pc�� L_���feÂސRBߐ<p>X�MC_ED'@�  H�Ni M�bG���MY19F�0EaS�L30� x �$OVSL�SDIsPDEXǓ�f֓$Hq�bV+��eN�a
���Pp�cwx�bw��=�c_SET�0�� @�Cr�%9�R)I�A3�
Vv_��bw�{qnq0-!�@� ��4BT� àAT�US�$TRCpA�@PB�sBTM�w�qI�Q�d4F��s�`.0� D%0E�P�b�rr�E1"�qQpd��qEXE�p���a��"��tKs�Rp&0�pU�P�01�$Q `X�NN�w���d���y ��PG|5� $SUB�q�%xq��q|sJMPWAI2$�Ps��LO ��1�
 �E$RCVFAIL_C@1�PÁR%P�0�#���Ȕ� ��
�R_PL|sD�BTBá���PBW�D��0UM��I�G�Q `�,�TNL ��b�ReQ�2���qP��@EǓ��֒���DEFSP� �� L%0� ��_8���CƓUNI�S�w�Đe�R)��+�_L�
 P�q"@��H_P�K�5��2RETR�IE|s�2�R���F�I�2� � $��@� 2��0D�BGLV�LOG�SIZ�C� ���Ud�"|�D?�g�_T:�ʥ!M�@C
 #EM⌭R��y0�8CHE3CKS�B�Po01���0.�0R!LbN�MKET��@�3r�PV�1� h�`ARp� �1)P�2>��S�@OR|sFORgMAT�L�CO�`�q����$Z��UX8�P!r�qPLIG�1ߛ  ˣSW�Im 6���,�G�AL?_ � $`@R��B�a��CS2D�Q�$E1��J3�DƸ� T�`PD�CK�`�!LbCO_J3����T1׿6� �˰C_Q�`� � ��PA�Y��S2u�_1|�2|�ȰJ3�ИˈŬƼ��tQTIA4��5:��6S2MOMK@�à��������y0B׀A�D��������PU��NR��C���C������4�` I$PIN�u�41�ž� ��:q�R~ȇ��ٯ� �:�h��a�֬��ց��1�'1R\uSPEED G��0�؅�� 7浔؅�%P7�m�F�p�U��؅SAM �=G��7��؅MOV	B� e0�� ��c2 ��v��浐�� ���c2@nPsR����İ$QH���IN8�İ��?�[��6�؂A���X����G�AMM�q�4$GGET1R@�SDe�zmB
�LIBR[��y�I�7$HI�0_�5a@c2E`@#A@ 1LW^U�@	�1a¬&o�ʱC�=�n S`�p �I_��pPmDòv� ñ'����mD��	ȳ� �$�� �1��0IzpR� D`T#|"c���~ LE^1�41�qwa�?�|�M�SWFL�MȰSCRk�7�0��Ѻpv���Z 0�P�@�9@���2�cS_SAVE_Dkd%]�NOe�C�q^�f�  ��uϟ�}ɕQ��}��Ѐ}*m+��9��ժ(��D �@���������b3 1�RA�Mam�7
5�#���^���Mtա � �YL��
A'�VAS	BtRna`7GP �B
Bl3
A%`�GSB1W? �2�2cЬ3doBB1M&@�;CL�8����G�b�1v���M!Lr� �N�X0�d$W @�ej@b��  @=�BD�BK�B� -�> �P����ycİ%X �OL�ñZ�E����uԣ ��OM�R/d/v/�/�/p��A�jM`���:e�_��� |��H  ��jV��yV��yP��ȗW�V��E��� Q�@pLT������NTP=��PMpQ}U�� � 8Tp�QCOU,�QT�HQ�HOY2`HY�Sa�ES��aUE� `"#�O���  b �P�0�rUN�pʌ3��O$�J0� �P�p^e������O�GRA�qk22�O��d^eITm�aB`INFOI1���k�a�k2��OI�b� =(!SLEQ(��a���`�foaS� ���� 4TpENAB|LBbpPTION|s�����Yw��1sGCF:��O�$J�ñfb���R�x!�]|ot�OS_EDŀNJ0� �N��@K��j��ES NU�w��xAUT,!�uCO�PY�����v�8 M�N���PRU�T�� �N�pOU���$Gcbn�l�R�GADJI1�2�X_B0ݒ$ ����@
��W��P�����@�l����EX�YCLB�IQRGNS6u��N0�LGO�A�NYQ_FREQZ��W���+�p�\cLA�m"����Ì�uCR1E  c� IF�ѝc�NA��%i�_G>mSTATUQPmMAIL�� 1���yd����!��EL;EM�� �7 DxFEASIGq2�� v��q!�er$�  I�`�"��ae�|&I�ABUq�E�`D�9V֑a�BAS��b�� [�Ub�r % �$y���RMS_TRC�ñj���Ca��`ϑ��,r���C�YP�	 � 2�  g�DU�����Ԣ�0�-�1��1���qDO�U�ceNrs��PR�30;p�rGRID��aUsBARS(�T�YHs$��OTO��I1��P`_��!�ƀ��l�O�@7t� � �`�@PORp�cճ��ֲSRV��Y)���DI. T��@�!��+��+�4)�U5)�6)�7)�8�҄�F��:q�M`$VALU|�%�ޡ|��7t�� Cu�'!�a���� (gpAN#��R�p0� 1TOTAL��[���PW�It�&�REGGEN$�9��SX��`sc0��Q���PTR��Z�$�_S ��9дsAV���t���rb�E���x�a�"^b�p��V_�H��DA�C����S�_Y4!�B<�S�A�R�@2� f�IG_SEc���˕_b`��C_����w���?r��%�b�H�SL)G#�I1��p"=����4��S�2̔D�E�U!Tf.p��T�E�@���� !�a����Jv�,"��IL_MK��z�н@TQ�P�a����2VF�CT�P���^�mMu�V1t�V1��U2��2��3��3��4��4����С����1�"IN	V�IB@N�; �!B2�>2J3>3J4>4JI05���"����p�MC_F,`3 � L!!�r�M= I��M�� [PR�� K�EEP_HNADED�!f�C�A���!����"O �Q I����"��?�."REM9!�Pϲ^uzU��e!�HPWD  �SBMSKG��a	!B2B�
#COLLAB�!��2������o��`IT���A`��D� ,�pFLI@��$SSYN� ;,M�@C>���%�UP_DLYzI1�MbDELAm �ј�Y�PAD�A��QQSKIPE5�� ��``On@NT�1� P_``�b�' �`�B]0�'���)3��) ��)O��*\��*i��*�v��*���*9�JS2R‎��?sX��T%�|1�{2ܐ�p|1�a���RDC!FW� ��pR�sR�PM�'R^��:b�2��RGE�p2��3d�F�LG�Q�J�t�SP9C�c�UM_|0��_2TH2NP�F@~o0 1� �0�EF�p11��� �l[P�E-Ds#AT Wo�[�w�B�`�d�A �p3�BfcAHnP�B+ ^E2gB�mOO��O�O�O�O�G3gB�O�O_ _2_D_�G4gB�g_y_�_�_�_�_W E_D5gB��_@�_oo,o>o�G6gB�aoso�o�o�o�o�G7gB��o�o&8�G8gB�[m�����ES����B\@ǡ`CN�@�1ZvE��^� @�o��m�IO�ፉIx���^APOWE!�� W�: �1�j�� �5%Ȃ$DSB;���֒ �h yCL@��S232s�'� ��0�u.���ICEU{���PE|V@��PARIT��Κ�OPB ��FLOW�TR2�҆�]���CUN�M�U�XTA���INT�ERFAC3�fUn��	�CH�� t� � ˠE�A3$����OM��A�0נI���/�A$�TN���Tо 8��ߓ��EFA� �8"!�Ґ�� u!��� O�� &*��� �����  2�� �S�0�`П	� �$3@}%�:B�Ŏ��_���D;SP��JOG��V�fh�_P�!s�ONq0�%�0���K��_McIR���w�MT7��AP)�w�>@"����;AS������;APG7�BRKH����G ��µ! ^���i���P���Ҏ���BSOCd��wN���16��SVGDE_OP�%�FSPD_OV%R�u �Dвӣ�OR޷�pN��߶F�_�����OV��SF�<��
�F0����oUFRAF�TOd��LCHk"%�OVϴ ��W[ ���8��Ң�͠;�  @� BTIN����$�OFS��CK��WD���������r����TR��T�_FyD� �MB_C 
�B��B����(�.Ѻ�SVe��琄�d}#�G)�<�AM���B_��jթ�_M�@�~��ቂ��T$C�A����De���HcBK�����IO�q�թ���PPA�ڀ������Տթ���DVC_DB��?��� �A��,�X� b��X�3`���3�0�����ϱU󳠈�CAB��0��ˠ��c� �O�w�UX��SUBCPU�ˠS�0�0� R����!�A�R�ł�!?$HW_Cg@A��!��F��!�p� � '�$U r�l�e�ATTRI��y�ˠgCYC����CA���FLT �����ث��ALP׫CH�K�_SCT��F�_e�F_o����FqS�J�j�CHA�1���9I�s�8RSD�_!聂��恩�_T`g�7�� �i�EM,���0Mf�T&� @�x&�#�DIAG��?RAILACN���M�0�"��1���XL��{�PRB�S  � ��C4�&�	^��FUNC�"��'RIN�0 "$�7Lh�� S_��(@���`�0��`A��CBL� u�A����DAp�a���LDܐð�����j��TI%���@�$CE_RIYAA��AF�P=��>#��D%T2� C���a�;�OIp��D�F_Lc�X��@�L�ML�FA��HRD�YO���RG�H�Z 7����%MUL�SE� �����k�$JۺJ����F�AN_ALMLV��1WRN5HA�RDr��Fk2$?SHADOW|�Ma���O2s�0N�r�J�_,}���AU- R+�?TO_SBR���3����:e�6�?�3MPINF@{��4���3REG�N1DG��6CV��s
�FL�W��m�DAL_�N�:�����q�h	����a�U�$�g$Y_Bґ u�|_�z��� �/��EGe���ð�AAR������2�G�<�wAXE��ROB��7RED��WR��c�_�M��SY`��Ae�:VSWWRI���FE�STՀ����d��EEg�)��D-�{2B��BUP��\V��D�ЗOTO�1)���ARY���R���Bbנ�FIE���$LI�NK�!GTH�R&�T_RS���E�N�QXYZ��Z5�V'OFF���R�R�X&�OB��,8d����9cFI��Rg��h􃻴,��_J$��F�貿S��q0kTu[6@��1�w �a�"�bCԀ�+�DU�¤F7�TUR0X#�e�Q�21X$P�ЩgFL�Pd� ��@p�UXZ8����� 1�)�KʠM��F9���ӓ�ORQ���fZW3	0�B�OPd�,��tp����A�tOVE�qeBM���q^C�udC�u jB�v�wL�wg��tAN=�Q�qD!fA�q ��=�}��q�u�q���0dC��"���ERϡj�	�E��T�ńAs�@�UeX��W����AX��F���� N�R��+��!+��  *�`*��`*��`*�Rp*�xp*�1�p*�� '� � 7�� G�� W�� g� � w�� ��� ��� ���đ��DEBU=��$8D3�h����RA!B������sV��<� 
��i�fA��-� ���������a���a ���a��Rq��xqJ$�`�D"�R9cLABOb8�u9�F�GRO��b=<��B_���AT �I`�0`����u���1��ANDfp�ຄ���U���1ٷ ���0�Q`������PNT$0~M�SERVE�Ny@� $%`dAu�!9�PO��[0���P@�o@*�c�x@��  $]�TREQ�2
\��Bf��j��D"2�{�" � _ �� l"T�c6ESRRub�I��VO`�Z���TOQY�V�L��@)�1R�Ƅ G;�%��Q�2E\�T0e�ף ,7�ř��]�R�A#� 2� d�@����r� �Y@$�p�t ��[�OC�f�� � ��COUN�TUQj�o@FZN_wCFGe�� 4B�F��Tf4;�~�\� ��
�ӭ�uC� ���M: �"fA��U��q: �FA1 d�?&�X�@=����eB�A<�����AP��o@HE�L@��� }5�`B_BAS�3�RSRF �CSHg�!��1
ש�2��U3��4��5��6���7��8
ל�ROO0�йP�PNLdA�c�ABH�� ��ACK���INn�T��GB$�Uq0� +\�_PUX��@0��OUJ�PH�H���, u��TPFWD_KAR��L@��REGĨ P�P��]QUEJRO �p�`2r>0o1I0������P����6�QSE�M��O��� A�S�TYk�SO: �4D�Iw�E���r!_�TM7CMANRQܨ�PEND�t$�KEYSWITCaH���� HE�`�BEATMW3PE��@LE��]|� U���F>��S�DO/_HOMB O>�_�EF��PR>a9B�ABPx�CO�!��#яOV_M�b[0# I�OCM�d'eQ��ZЊ�HKxA� �D�QG��Ue2M������cFORC.CWAR�"�ъ��OM�@ � @�r�:#�0UHSP�@1*&2&&3&&4�A��*s�O��L"�,�HOUNLO��c4j$�EDt1  �S�NPX_AS���� 0+@ @��W1$�SIZ�1$VA����MULTIP�L��#! A!� � $��� N$S`�BS�ӂAC���&OFRIF�n�S���)R� NF�ODBU$P���%B3=9GŸ�Ҫ�y@� x��S�I��TE3s�r�cSKGL�1T�R$p&���3a�P�0STMTd1q�3P�@5VBW�p��4SHOW�5���SV��_G��� Rp$PCi�oз��kFB�PHSP' 1Av�Eo@VD�0vC��� ���A00޴RB% ZG/ ZG9 �ZGC ZG5XI6XI7�XI8XI9XIAXIB�XI ZG3�[F8PZGFPXH��XdI1qI1~IU1�I1�I1�I1�IU1�I1�I1�I1�IU1�I1 Y1Y1YU2WI2dI2qI2~I2�I2�I�`�X�IQpT�X�I2�I2�I2�I2 Y2Y2Y�p�h�dI3qI3~I3�I3��I3�I3�I3�I3��I3�I3�I3�I3� Y3Y3Y4WI4�dI4qI4~I4�I4��I4�I4�I4�I4��I4�I4�I4�I4� Y4Y4Y5�y5�dI5qI5~I5�I5��I5�I5�I5�I5��I5�I5�I5�I5� Y5Y5Y6�y6�dI6qI6~I6�I6��I6�I6�I6�I6��I6�I6�I6�I6� Y6Y6Y7�y7�dI7qI7~I7�I7��I7�I7�I7�I7��I7�I7�I7�I7� Y7Y7T�VPz� Uc�� l�Dנ��
>A820��5��RCM2����MT�R��|���Q_��R-��ń����[��YSL�1�� � �%^2��-4�'4�-Y�BVALU��Ձ���)���FJ�IgD_L���HI��9I��LE_���f��$OE�SAbѿ� h 7�V?E_BLCK�|�1'�D_CPU7� � 7ɝ �����E����R � � �PW��>�E ��LA�1Saѝî���RUN_FLG�� ������� ��������B��H���Ч�ɠ�TBC2��� � _ B��� br�p W?�eTDC�����X��3f�S�T!He�����R>�k�?ESERVEX�Ԅe��3�2 �d��� �X -$��LENX��e�Ѕ��RA��3�LOW_�7�d�1��Ҵ2 �MIO/�s%S80t�I���"�ޱH����]�DE<m�41LACE�2��CCr#"�_MA�� l��|��TCV����|�T�������@0Bk�)A�|�)AJ��%EM7���J��B@k�)X�|���2p �0�:@q�j��JK��V�KX�����ы�J�0����JJ��JJ��AAL����������4��5�Ӵ N1��� ����LF�_d�1� � �CF�"�� `�GROUP���1�AN6�C�#~\ REQUIR�Ҏ4EBU�#��8�$Tm�2���|�ё %�� \�A�PPR� CA�
�$OPEN�CLOS<�Sv��	k�
��&� �<�M�hЫ���v"/_MG�9CD@�C ���DBRKBNOL�DB�0RTMO_�7ӈr3J��P ��������������6��1�@ ��;$���# � ���'��-#PATH)'B!8# B!�>#� � �@�1�SCA���8I�N��UCL�]1� C2@UM�(Y"��#�"������*���*��� P�AYLOA�J2=LڠR_AN`�3�L��9
1�)1CR?_F2LSHi2D4LO4�!H7�#V7�#ACRL_�%�0ȑ'�$��H���$yHC�2FLEX�u;J#�� P��4�F߭߿���0��� :����|�HG�_D����|���'�F1_A�E�G6�H�Z�l�~���BE������ ������*��X�T,� C���@�XK�]�o�^Av�T&g�QX>�?�� 4TX���eoX������ ������������	t-	�J@� �/�`M_q~�۠AT�F�6�ELHPѬs��J� � JEoC3TR�!�ATN���v�|HAND_VB���1��$� $�:`F2Cx���S�W�A�"�� $$M,00�_�Y�ni��P\����A@��� 3����<AM��_AmA|��NTP�_DmD|P\ G��E�STaM�nM�NDY��� C ����0��>7_A>7Y1@�'��d�@i`�P� ������"Qs$�� O�4D'"��xJ���ASYMl%A�� l&��@�-Y1�/_�}8� �$���@ ��/�/�/�/3J	<��:;�1�:9�D_V�I�x���V_�UNI�ӝ��cF1J ����䕶�Y<��p5Ǵ �y=6��9��?�?>��wc�4�3���$� ASS  o���s�  ��{�h�VERSIO�Np�~��=
��IRTU<�q����AAVM_WR�K 2 ��� 0  G�5z�������&� 9 �	8�)�L�{����:�w�^�|�(ܛݧ�7ѭ�����|����BSPOS�� 1��� <��A�S�e�w� ������������ �+�=�O�a�s����� ����������' 9K]o���� ����#5G Yk}����� ��//1/C/U/�>��AXLMT��X#��%�  dj$I�Ns/�!i$PRE_EXE�(� �&)0�q�������LAR�MRECOV ��ɥ"
�LMDG� ����[/LM_IF �� �!X/c?u?�?�?�:Q?��?�?�? OM, 
0�8O�4�cOuO�O��O�NGTOL � ���A   ��O�K��PP)�O ; ?6_,_>_P_{� $BR_�_ w�o_�_�_�_�_�_o@�_'oo7o]o�!��O �o�o�o�o�o�o�o�+=Oa�PP�LICAT��?��� �J`�Handling�Tool �u �
V8.30P/�33�@lt��?
88340�slu

F0�q��z{�
2026��tlu��_�7DC3�p�J  �sNone�lx� FRA������B��TIV�%�s�#~��UTOMOD� �E�)P_CHGAPON������Ҁ�OUPLED 1��� ��"��4�uz_CUREQ7 1��  � >�>�*ސ�4��!���x�~� ��u��Hm����HTTHKY�� ��w���7����%�C� I�[�m��������ǯ ٯ3����!�?�E�W� i�{�������ÿտ/� ����;�A�S�e�w� �ϛϭϿ���+���� �7�=�O�a�s߅ߗ� �߻���'�����3� 9�K�]�o����� ��#������/�5�G� Y�k�}��������� ����+1CUg y������ 	'-?Qcu� ���/��/#/ )/;/M/_/q/�/�/�/ �/?�/�/??%?7?�I?[?m??��P�TO��@����DO_CL�EAN܏��CNMw  �K >��aOsO�O�O�OD�DS�PDRYRO̅H	I��=M@NO_'_9_ K_]_o_�_�_�_�_�_8�_�_J�MAX�p�4�1���aX�4"��|"���PLUGG����7���PRC�@B�;@?K_�_ebOxjb�O��SEGFӀK�o�g�a;OMO'�9K]�o�aLAP �O~Ǔ����� ��/�A�S�e�w���>΃TOTAL-fVi�΃USENU�`��� ��䏺�P�RGDISPMMC�`e{qC�aa@@}r���O�@f�e��_�STRING 1�	ˋ
�M�ĀS��
`�_I�TEM1j�  n ����������Ο��� ��(�:�L�^�p����������ʯܯI�/O SIGNA�Ld�Tryout Modek��Inp�Sim�ulatedo��Out.�OV�ERR�@ = 1�00n�In c�ycl"�o�Prog Abor8��o��Statu�sm�	Heart�beati�MH� Faul����Aler���ݿ�π�%�7�I�[�m�� �3f��1x����� ������*�<�N�`� r߄ߖߨߺ�������8���WOR�`f� L���&�t����� ��������(�:�L��^�p�����������POd�����d��� %7I[m�� �����!3pEWi��DEV�� ������/ /'/9/K/]/o/�/�/��/�/�/�/�/�/?PALT��81d�? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnOp�O�O�O&?GRI` f��AP?�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHo�OR�̀a�OZo�o�o �o�o�o&8J \n������<�noPREG<>%� �o�L�^�p������� ��ʏ܏� ��$�6��H�Z�l�~�����$�ARG_L�D ?�	���ӑ��  	�$�	[�]�����ƐSBN�_CONFIG S
ӛ&�%� ��CII_SAVE  �E�<�Ɛ�TCELLSET�UP Ӛ%  OME_IO���%MOV_H8������REP�l����UTOBACK�t�0�FRA;:\� ����_�'`���=�{� J� 	� �����ͿĿֿ�6����	�1�C�U�g� yϋ��Ϸ������� ��ߜ�5�G�Y�k�}� �ߡ�,���������� ��C�U�g�y���\��a�  )�_��_\ATBCKC�TL.TMP DATE.D;<��	�p�-�?��INI;0�p�8��MESSAGT�^�_�ېi�ODE_D��W�8��H���O����PA�US��!�ӛ ((O֒��
�� *N<r`�� �����"��~��TSK  ��x=�C�	�UPDT���\�d���XWZD_ENB\�4���STA[�ӑ�őX�IS&�UNT 2�ӕ`� � 	 S
/��2//V/A/�z/e/�/�/�/�/�M[ET�`2�P�/�?�/<?�)SCRD�CFG 1C�`��\�\� 1?�?�?�?�?�?�?6��QX��??OQOcOuO �O�O O�O$O�O�O_�_)_;_�O�O���G�R����zS��NA���қ	�wV_�EDZ�1e9� �
 �%-��EDT-h_ʪ�_o�`/^���-��_��	������_�o  ���e2�oɫko �o�6k�o!hozo�o�c3Y�o��o�n���4F�j�c4 %��r���nN��� ����6��c5�a�>� ���n���̏ޏt���c6��-�
�Q��n�@Q�����@�Ο�c7�� ��֯��n���d�v�����c8U��_����0
 }~��0�B�ؿ�f��c9!ϑ�nϵ�  }Jϵ���Ϥ�2φaCR�oį9�K���߀�����n���zP�PN�O_DEL�_xRGE_UNUSE�_�vTIGALLOW� 1�Y~�(�*SYSTEM�* 3	$SERV_GR�R 69���7REGB�$d� <�9�NUMg��z��PMU�� 5L�AY�  <P�MPAL[��CY'C10����������ULSU��{������D�L�N�BO�XORIk�CUR�_;�z�PMCNmV��;�10��>��T4DLI�4�V���ߨ���'9K]oR�zPL�AL_OUT �Dcc�QWD_A�BOR��	��IT_R_RTN���Y�� NONS8�� �CE_RIA�_I��<FF_1�4e :[�_PARAMGPw 1�w�`_����Cp�  .� � �� � � � �� � � � �� � �  D�X $3!g-�<$��H$�T$� D*X � X "� B�kD1� 9X @� 6�?� <HE��ON�FIy���!G_Pv��1� �e �U??0?B?T?f?x?|�?�!KPAUSX�s1�UR ,Z� �?�?�?�?�?OOO TO>OxObO�O�O�O�OмO�O_�2O_�ey�PCOLLECT__�Y[ 4cGWEN��I�"cR Q�NDEOS�W���1234567890�W�S�p5b�_�Vy
 H�y)�_#oS��_oho T�AoSo�owo�o�o�o �o�o�o<+� Oas����� ���\�'�9�K����o��VQ�2W[ �� 9W�VIO �YcQyH&�8�J�l\��TR�2؍�(��
��j�� � ����%�_MOR҂!� + �'� 	 �5�#�Y�@G�}�k����Ӂ"��2?�!�!3 ҡ��Kڤ��$R_#�*_	�:Q:RC4  �AS yC  x�=A3!z  BC!�P�B/!�PC  @�*����:d��
�IPS$����T��FPROG %�*6߼�8���I����&RҴKEY_TBL  )V�R:P �	
��� !"#�$%&'()*+�,-./�W:;<=>?@ABC���GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~�������������������������������������������������������������������������������������������������������������������������������������������1��L�CKۼ3���STyA�д_AUT���O(��U�INDxtTD�FQR_T1_�Q�T2��7$����XC� 2����P�8
SONY �XC-56�9Q}����@���u�} ��А�HR5��cT0�B�7<T�f�Affrꬿ���� �������5� G�"�k�}�X��������������ǼTR�L��LETEG���T_SCREE�N �*k�csc:U$MM�ENU 1&�)  <��� y��Ã�= &sJ\��� ����'/�/]/ 4/F/l/�/|/�/�/�/ �/?�/�/ ?Y?0?B? �?f?x?�?�?�?�?O �?�?COO,OyOPObO �O�O�O�O�O�O�O-_ __<_u_L_^_�_�_ �_�_�_�_�_)o oo _o6oHo�olo~o�o�o �o�o�o�oI 2�X�hz���� _?MANUAL�ߕ��DB��L+�DB�G_ERRL��9'�� �\��n����NUML+IMK�d �p��DBPXWORK 1(�I�ޏ�����&�ŽDBTB_@ )��������qDB_A�WAY�_�GC;P  �=�װ�~��_AL��D�z��Y���M � �_)� 1�*����
�͏����6�@�_M&{�ISAЉ�@B�P��ONTIMJ�& ��p�ƙ
�ۓMOTNEND߿�ڔRECORD ;10}� �>�?�G�O����?��� 2�D�V�h���p���� ��*�߿�Ϛ���9� ��]�̿�ϓϥϷ�R� ��J���n�#�5�G�Y� ��}��ϡ�������� ��j���C��g�y� ������0���T�	� �-�?���c���\��� ��������P����� ;��_q����� (�L%�4 [�����^ t�l!/�E/W/i/ {//�//�/2/�/�/�??�/z�TOLEoRENC��B�ВL���CSS�_CNSTCY ;116�  ?Β�?�?�?�?�?�?�? OO&O8OJO`OnO�O��O�O�O�O�Oc4DEVICE 126� b�*_?_Q_c_ u_�_�_�_�_�_�_?��d3HNDGD �36�Cz�^LS 24]�__oqo��o�o�o�o�o�_e2PARAM 5��B��t�dc4SLA�VE 66�e_?CFG 7��gdMC:\e0�L%04d.CS�V�o��c|�r�"AM �sCH�p&a&�P�n��w��f�r�����ÀJP��>��\_CRC_�OUT 8U�����oEpSGN �9U�Ƣ��\��12-OCT-�22 17:27ܬp�0��4:�41�p9V UBu1�݁�nހ���o��Im��P��uG��@uVE�RSION ���V3.5.�11E�EFLOG�IC 1:ݫ 	6��|�C����^�PROG_EN�B����͢��ULS�{� ��^�_AC�CLIM|���Xs��WRST�JN[���ţ�^�M�O��¡Zr,�INI�T ;ݪs5� �*�OPT$p ?�	i�B�
 	�R575�c��74j��6��7��50��R�Ƣ2��6��X�y�TO  ���?��Y�VP�DEX�d����@W�PATHw A��A\E������7;IAG_G�RP 2@�k�,�"	 E� � F?h Fx� E?`�D��@û��V1"�ü��T0�K�9�Cf�py�pY��dC�pq��B�i�ùm�p4m5 7890123456���;����  A��ffA�=qA�ةpхA��WHAĩp������?�A��Mk���@��tp�p��W0�A�T0T0�pB4�ü Qô���
����(�A�A��
=A�L����A��
A�Q��A�������� e�����e� Pe�:�_�{A�d������dѩp�������A����������r߄ߖߨߺ�@�EG��A@�p:�RAU5d�/��)��#P�d�l������"��4�F�@�Pz�AJ���c�?��9p�A�3\)A,��A&����0���������@�cP�]���AW�P�J��C���<d�4�-d�%G��(�:�L�^�@� ��$HZ��. |����bt�  2Vh�xm� ����[���s������=�
==�G���>�Ĝ��7���8��b��7�7�%�@�;�\"&�p�.%���@�Ah�p9 A���<i��<xn�;=R�=s���=x<�=�~�Z�;��%<�'�'�~ �?+�ƨC�  <(��U� 4"�;���&����%ùf��@?Œ?�? @?R?g��$^?�?"?�?�?�?�?�?�?)7�L?S�FB$��/"Eͽ�>OG��ΐԬq��sD�L4�x�CA��Gb�t� ����-_7_�C��_�;�/_�NED  �E�  Eh� 	D[PbRD_¿�_�86��_�_
z{_�_w_o�K:o@bù Qm)o�o�oo�o�o�o��o ɼCT_CO�NFIG ���Yt؃e�g��ԱSTBF_TTS�
ęVs3����
�iv[�MAU����Y�MSW_C5F*pB�  �Q��OCVIEW}pC�}����_�!� 3�E�W�i�;������ ��ȏڏ�{��"�4� F�X�j���������ğ ֟������0�B�T� f�x��������ү� �����,�>�P�b�t� �������ο��� ��(�:�L�^�pς��|KRC�sDJ�r!� �κ�������7�&��[�otSBL_FA?ULT E���x>u�GPMSK_w���pTDIAG �F.y�q�IU�D1: 6789?012345��;x�MP�o!�3�E�W�i� {������������`��/�A��X W!��J�"
��vTR'ECP����
���� �M�(:L^ p�������  $6]�o�l���UMP_OPTIcON_p�ގTR�rt`s���PME^u��Y_TEMP � È�3B��pp �A  �UN�I�pau!�vYN_?BRK G�y���EMGDI_STaA%�1!G%NCS#1H�{ �K��9�/_}dd�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO��O�O�O�O �I�!�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo �JO�o�o�o�o�O�o �o+=Oas �������� �'�9�K�]�wo���� �����oۏ����#� 5�G�Y�k�}������� şן�����1�C� U�o�]�������ɏ�� ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�g�y��� �ϧ�]�ӯ������ %�7�I�[�m�ߑߣ� �����������!�3� E�_�q�{������ ��������/�A�S� e�w������������� ��+=Oi�s �������� '9K]o�� ������/#/ 5/G/ak/}/�/�/� �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OY/KO uO�O�O�/�/�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oQOcOmoo�o�o �O�o�o�o�o!3 EWi{���� �����/��o[o e�w������o��я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�S�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�K� 9�g�yϋϥ������� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�C�U�_�q�� 9�Ϲ��������� %�7�I�[�m������ ����������!;� M�Wi{���� ���/AS ew������ �//+/EO/a/s/ �/��/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O =/GOYOkO}O�/�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo5O'oQoco uo�O�O�o�o�o�o�o );M_q� �������� -o?oI�[�m���o�� ��Ǐُ����!�3� E�W�i�{�������ß ՟������7�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �/�9�K�]�oω��� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ���������'��C� U�g��w������� ����	��-�?�Q�c� u��������������� �1�;M_�� ������ %7I[m�� �����)3/ E/W/i/��/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?O!/+O=OOOaO{/ �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_O#o 5oGoYosOeo�o�o�o �o�o�o�o1C Ugy����� ��o�-�?�Q�ko }o��������Ϗ�� ��)�;�M�_�q��� ������˟ݟ�	�� %�7�I�[�u������ ��ǯٯ����!�3� E�W�i�{�������ÿ տ�a���/�A�S� m�wωϛϭϿ����� ����+�=�O�a�s� �ߗߩ߻�������� �'�9�K�e�o��� ������������#� 5�G�Y�k�}������� ���������1C ]�Sy����� ��	-?Qc u��������� �$ENETM�ODE 1I^��  
  (/:+
 �RROR_PRO/G %*%}/��)X%TABLE  +h�/�/�/��'X"SEV_NU�M &"  ��!!0X!_AU�TO_ENB  qD%#U$_NO21� J+9!2�  *�u0�u0�u0�u0(0+t0�?�?�?N4HIS3
 �G;_ALM 1K.+ �u< +�?/OAOSOeOwO�O�?_2T0  �+s1:"�J
 TC�P_VER !�*!u/�O$EXTLOG_REQ�6s�E9 SSIZ)_�TSTKFYc5��RTOL  �
Dz�2�A T_BWD�@�P<6ܯQ8W_DI�Q L^G48$
?"�VSTEP�_�_
 >�POP_DOh_!�FDR_GRP s1M)B1d 	�O�fo: W`�������glp�w�qŗ��I ����f Wc�o�m�o�o�o�o (L7I�m���zA�f�A�؟�>�Β� 
 E��	�q� @(�C��<�'�`�K��C`}dC��N���B�{��F�@7UUT��UTF�Ϗ�j��s���sOHc�EP]��O���#M��*�KA�����?�pF��:6:N�r�9-�z���c ����������+FEATUROE N^�P>!�Handl�ingTool �� mpBo�English �Dictiona�ry�
PR�4D Stڐa�rd�  ox,� Analo�g I/O�  �ct\b+�gle� Shift� � !*�uto S�oftware �Update  �fd -c�mat�ic Backu�p�IF O���ground �Editސ�g �R6Came�ra3�F7�Par�t��nrRndIym���pshi���ommon ca�lib U���n�����Monito�r�CalM�t�r�Reliab�L��RINT�Data Acq�uis�Z�ϠC�iagnos��0�<��almC�ocum�ent View�e�\���C�ual� Check S�afety��  �- B�Enhan�ced Us��Fyr���8 R5��xt. DIO 6�fin� (�@ϲwend��Err�=Lm� D p^��Z��s	�EN�r.��հ �P�rds�FCTN MeKnu��v8���m��FTP In'�f�acN�=�G��p �Mask Exc���gǱisp��H�T^�Proxy �Sv��  VLO�Aאigh-Sp�e��Skiݤ e�f.>�Hf�ٰmm�unic��ons��
!
��ur�E�'�7�rt F�4�a�conne�ct 2;�Inc=r`�stru����� SpKAR�EL Cmd. �L��ua��OAD�*�=�Run-TiNưEnv� �D;�^(�el +��s���S/W�.{�License���
����ogBo�ok(Syste�m)蔭�JM�ACROs,��/�OffseS�Z�M�Hٰp��� j73�ΰMMR��l�3�5.f��echS�top��t�R� 7ize*�Mi��O� 2�7�x��0���n�miz��odM�witch����a�.�� v���O7ptm��49����fil��ORD���0�g�� 849~6�ulti-T�������CPC�M fun,��.sv�oO����� �^�5�Regiҷ�r��	�!2�ri���F�  H59�k�1�Num Se�l*�  74 H|��İ Adju����adin��O� y,[���tatub��\У�������R�DM Robot���scove� ��d em(�ٱn�� SW��Servoٰs�ꒄ�?SNPX b���1��g P�Libr<���1�ڐq 9� ɰ.30g �o��tE�ssag�� f��@ �e����"g��/I�_�
�I�TMIL�IB���� P Firmn���^�FAcc����0���T�PTX���510.� eln�����x����H573��rquM�imul�a��� 2�ToMuz�Paxѩ1� �T��6���&��ev�.��IUSBg po����iP�}a�� 0\sy nexcept��|3 <� \h51 �����oduV #��9��Q�VN�k"6PCVL{&�^�}$SP CSUI��d���+XC��a�uҠWeb Pl���t? �#S��\" 	2�������S�&ުz�V?8Gridplay��&� ���8�-iRb".� �@ � R-2000�iC/165¦ �d+�+�larm �Cause/1 e�d�<0:�Asciyi����Load��V4�3Upl�0�_�CycL�c�m�or�i����FRA[�a�m�) tdt��NgRTLi�3Onݐ�e Helݨ 5�42*�PC`ρ�4��`�]�1trߵ4�8��ROS Et�hv�t[���10�\ҠiR}$2D ;PkߵDER>1�E����of�A��ΰ�FIm��F�� z���64MB DRA�Mު�@:�9RFRO<A[�Cell3� �����shrQ
��ZcЛ��ÍUk�p� p�ide�WtyL�sL��|0\z�!Ctd���.��@"EmaiF��li���+�\��� R0�qZ$Gig�E�N�4OL�@Sup"��b�W3oa�~�cro������4���QM��Fauesat�A>�j�� miH9.dVirt��W��0{&ImM�+T����}$Ko�l Buir��n�յ'APL�&4��MyV6� "�0�*�CGP�l���{RuG�'p�{SBUW��RQ�)K�&cm\ :��z��fX�)O�v�v�(TA�&spoҠ�-�B�&��
 I�\E �P�+�CB'fg-x��&"  �E��sv�b��vv�3���S_k��TO;-�E�H�f6.
�E�vf�x_z�)�V��tr >�)�hZ%.�F�&  � ��r���*�G�&�� �њr����H��Р^JzCTIAc�pw�4�LN�1�Mr�"C #[��g�"�M�$-�P2�~T�@�����vxui�-�SD�&�S�&�*4�W���2.pc�)VGF���fxwʪVP2AU \fx���N��if�u���"inVPB���)���s�D��*�a<�s�F�5 M��zs�I��c�{&�Traİ��U,p  ��<��2��<RDp	�N��HY�<��p��-��H����Øp)����y �ϭ����ħϞ��rд����í�4+���'9Ly���ӎ��yߞ9ӫ�c3�U���B�O�q�u�y�kߍӍSy*�ߞ��\Yy����k��W���ӄ�Yyx����:�	�ߞ�����5�o��e/�Q��,y�K�m��g�^~���us�2��A��������F�������y�)���|��<��1�m�.�+�M�Ϗ�8G�i�7n��c���1�� <����W������7�{����6��Z������uk<��[�|�!�3�?�ϔ��iB\�g���_��{�x@.��wrs�t���B�� H#68��@H)xT@J�EENDI?N��tql[}
_��w�P�TQ y(��I) "���PA���T�/��'85/A#bs;/ �C/U/�,q�/B�Gp`�/�#��/�"36��5�R ?!2epai?5!:/Y4W���%INTo?e?_.q�?�4)��?�2pa2g��?�F O�?A�a�d6?��t ZUD2�gunOOqC533�R?�D�0u�O�/�Mcam���OO�LNT� ?��P_�Ĕ�0_QR7�L_�Cfi._H?_,_�f'R50�_�SAF�-F�_�7�w.v�o��_�_8�/�dM� Cbo���o�bv9rEo��paa�oaDx�@�osF-AS"-sS�p'Is(�PC�esXPL�O�tlo�_�ut\a�Oh%a9fvh%- B��/�����C�$��sr�p�?@_�?`w�}�bA�����h�`��]T�<ˏ�sgch�o2s�t��CG\s;��u1s�?���Sg�/�gG J����GDǟri$"�o�gdiʏ�!�fd���?h%J364S��Tut�o�O �?s����F�_��� �E�0���D`!�)�`NO4E�O�i$II���iwjOl�ž��>�?*�lb
��V��vjr/��
���7���2��_�?zG7\2O�E G��Ϲ?���1� ޯ&��_d�oi�8��c��50�>�x�Ͻ�"L�o�h%����dj9��﴿ƿؿ�c� u9p9�C� j9{�E�2�L��Ek,B串 ����oS_e_�&/���O}�j94JϬ�duZ��U��=d;������8���r7�Dh�u���;]m AT��������f�a���M����P��-4r V��O"3 #S�dwc�P��in�`�a�?& �HTuRef���I
�?hc�g�r"���q.JG"�er�M/��/ �/LRA�^��uH71�/�tC9K�/<eTXP/?i�9k1/m5k.f��3riR�eHG�/ƪ/ cr�NHG�Rf?L�iY�7�hOuX��H\mO��oρ� ;H��DD@�O��*�<��:I�?�?��d�R�_ 3hd�ghgOO��_���gmh�_h�m ��XO�o|O�O�o�O\/$�o0�f�gm�o`���`e۠;iov���yt��"��uR60���#tmo_�3#1��fdr,�op7��_����lp�>oh��冬~� ߏ�dgts���&dޏ�/�o�o
��J?<�vrF���v.�R���Ɵpld�5�6�%4�0/���re�eK�m�XP)�KCO*O|%56?�OZ�` o~����E$io��0��jߠ���l ����3OR��LOFvod��_IF��$�� ߪ�dDߦX!B� Uce��ft�4 ���(M�O�5)e?Ƕ/���1?Q�D�uk�'�|� ���`�boto�����-���6�p�eS ��on*���^�lB'�����Տ_�q�_�rdk��4f��C(ҿȿ ¯ԯ������̟��𒜩��
I��5s71��t�adi3f9Tar��l�ofk0�������vPa�@�� PJ��|*`��������et�&4epg���ed��� E�5�RI � H552n� 747�21�p�WelR78��,� �0ETX�J614���ATUP  wwmfh 545�p��"6�pk�V�CAM  7\a�wCRI@ EwD" G UIF)�!28  j�C�NREM�`�63��a�SCH  �4C DOCV�� CSUi�!0� D sEIO�CE�54�#R�694 we!!ES�ET=S#!3!�a 7�3!fanuM�ASK��PRXY�_"7� �0�'OCO��"3=P[�<#"�ER J�" x7�!!J774#!;39�  Eq�G1��LCH 0#OP;LG%J5000#oMHCR)%PS�1.7#MCS 4D"�0�4 O#J55 [#MgDSWe!Y1MD#1�s#OP#1#MPR$07�0w"0�#�  Σ#PCMX �#R0 A�#� &�00�#� 0( �&0�$50( �#�PRS� 3J69\03FRD@ 02�RMCNy�ndM��93 SwNBAA�800�@�HLB  "Lo��SM�A0 (W�w"4 onit#!2�  II)�TC< [#TMILe �B��`0"K3�@TP�A� �QTXa�t�\j�@EL�BM25�0`0/D8��$78n�mon�195d vSD95\FUEC 0OP� UFR@ ��;!�C@ \�@;!O�0p�t"VIP�@#� I:�@0�!CSX� �#�WEB �#HTT. \stB24 �#�CG�Q#IG�Qtwopm�PPGS!�f�PRC�@SH7�$��w!6( �8��!�[�R RBB- Ci��B01rogw!#IF#"098-!!` ��@�A64�(AaN�VD�!Ld�1h 6a6�8( c�`d SR7^c!te.p� 0ka�ч@�bc`� CLI�$0?�sb$c9G MSp�"5a�` - A� wSTY�@al �@�CTO �CJNN�0J98�ORSp�0G��b�g J�`�OL�1Abn: S�ENDu�to�!L��Q���@*r#SLM�� 8�"FVR� M�CHN0CSW!SPcBVP�� PL� �ds �qV$0�cCC�G $p�aCR�0
�Np�QB� 87.f:�QK� j70*`�p��0'3CSqToo��CTQ���qTB$�P�N��@n;pq�C�@�Q#�� �p, #�p ��. %�$07#%�� `8D#TC� QSQ"TE� [#m� �tTE� gt"m�P�T�TF�Q[����@�#C�TG�Q�"���@�#C3TH `�TTI�@#�CT'Qeqs�PCTM�@SC�$0gS�^�0bodyqP�@�  ��� �1� d��q�a�us�a9��P[�qW4 `@06; GF `8��V@VP2@ 623�R i��@j?�g� `n��g�B `" g�D� `��g�FX mna�"PVPI��+ G V��!#V	`  23ƱRVK�@Np�@CV��Q31�934.��vo R�er�ne땗����i$��r���h��0�A���37� �<�"�\srv�����b�3b�- S�r�B"0���A�J�935땿B�5 (S�O���g ��1�1�R|�j9�3땷b��EN�5��� awm�SK� Lib��� ���������@	 �"|�h�h�#땼�b�wmsk�n�E����q���py&E�  ���!�0�2�t Fuïբ6xۯm��uji-�	I&���8k��8!�� ��땼P��2�2��2�Mai'�on@��_�/r�;pڦh;Ѐ;�G��_r���!��4�\ֶORC��+�5.�� "T¦TP��,hQ�652�1��4���<�xk�����ߦ�%t�P��QrֶSB�� ch_����)��t!0�B�"̿ h�h 땇�;���c������������>�Rp� �\toֶ3���cl�W��2p�"����� �����F����b@� Qt�a�϶0t��2ܐFsȒ�76�p䵝t	� Ad���5�82��ob�|*�{�\a��FMpQ ���A�migֶ�I�or�wI�.j�rfm��Fc����@1�EYE~� Iw���R���4�,K2Х70.�E��ld,�C�� 1�PTP]���.�"AD.�F�&3 k���ask��ȍ`4����۳dֶے��ER~�7 R�ƫ/�`T�?)�e�rv榀G?Y?k?}?�?�?ӹapa��	d����rƚ4�M��te����7H9!J�d/���G�p�ac�T��<6�b`�/� QO��$vc>�",@Vg����eYW�2�5/� BJ�h�F��R5:�d���0�`��@��I_�raj��e��he}�$`��e5(Xa�@��et���1Otdj��,�_�h�\	UI�/k�jAo�FO��`^���F��r��qW65q���K z�'6ڦus W'�Cb,'��'?��n��MFR��;]�lf�ǯ�fr>֛�w�p�/�,��_U[ǀ�мn�x'_i�{��� ��O���pJ���[@�o�in7L�O�9�\^ � 1R����+mi2״h� �j��҇- f�n�t >�MA H��I  Hw5529� (Cߑ�21��leR�78�c�ߒ0AcaJ614��~�0ATUP��ܓ��545�t-f�l�6yE=�VCA�M�tFLXC�RId���o�UIFnULX �28���mo�NREu'��6q3��WQ��SCH��=Cn�DOCV�gϠwCSU1�cxr��0$�;EIO�C%tx\c��54��oQ��9T�;�ES;ET�Temo?�S��/��7S�{�MAS�K��70��PRX�Y�T�`��7��`�O�ߐOCOe�\?�3�ô`>��0{�?���|�-��on G�?�39!'ߑõ H82LCHd���@IOPLG.�tCGM?�0��GО��MHCR�Go�S��/1_�CS4�cg�m��50T��?�5x$�[���MDSWMfb.�D�����OP��oX/2L_�PR���K�����{���88�3n�CM��0iAE,��0�Ő`~�5#�\h88�+�?��D���.?���4��0D�3��o�S4�����9��,iFR�Dd�/2E/��M;CN5�H93�K�oSNBA�U"R��7HLB��SM�՛�8��T���J52�Sa�ߐTC4�\�TTMILe��P��䴝A|�TPA���T�PTX��5��TE�L�ԫ�0䴈P��8`�˳���K�95��v��95��888��wUECd�rt �GUFRd�__�Cd�;2e-�VCO4��GVIP�;��I�T;AX~�CSX������WEB4����H�TT4�ka��2T�2�M/So�G#��Q�IG��< .�IP�GS=t\rxO�RC��aߐ7�/a��16D�s@>�R7#��! ��Oq�Ҥ��P��Ҷ�;�A���KÑ�$�0 �"��4����NVDx4���#�Adap���8D���68����R�7���P��D0��a��o�bܠ. CLIƔ�l\-C���CM�S�'��4�d "�ްSTY�[�CTmOT�tl��NN����ORS4�;�1 ��7ltiΰOLS�( AE���0�T���L��6�@���9@ ��L�M4�HV o�V�R���CS��shc>�PBV4䫁/��PL�
APV��u;st>�CCG4��0�nCR�4 H5���B���K�H573���?�����\cms�#�st.~TB���! �
�7�C�ԓ�?"�Oawsh?"��I04?"��3�TCd�K�\A 4�\sl"EĤpP��� 4�C[П"Ԥ�8c��"4�(��CT�F��c��"���C[TG�73m#G䖫THd�h� �Il��K�CTC�59m�'CTM�5M����Q0��re\g�P ���12��04��h���%S��13M�CTWd�9[@_�GmFd�SE]�P2d��t+��2�ա �2d�e[ll��PBd�I����1Dd��a�1F��t;ap VPId��ÓCV�!Vq��UA���CVK�ۣCV>#�coreL���H"�Hp!�HK"�H�atc�J�H�4$�I� �IL0H�I�2��H��H+2�IL�Y4p=�H���Ie\a�I�2 Z93�I{�H�@�NZ+��H 1��K48�Z<A�Ht{�Il �Z;"�O�Fs\!�Hk"�H {"@o�F[�PZo�Z���J��Tok�РH��H�\��Il�Z��Z2�=[ng-[gToo��I�p�j(�njrob9t_�Xbt.�JL� iur�o�I��i�!���F��POz�lin�g�j��y���Y"r�^zۢ�I�p��Gea�t^j�]��Z��_je �����_��lkҠHAm,��H|��Z��A�I�  �_�  ����Gvhm�J{�sqvnj���H49\�Jz�@L�Ij749{P�Zt\jNj�@_�"g.pjmcal��0�fu�J��^zh�m-��_bg���o�\rͫ �1�H! j���;����MT "�(�Cu�zk��bgft��JlpX���GCT�"���Gfc]�˝2�6\fߟ�926�l\� Ίu�>m��;�Mul?�Q��#7\^�K���7-[˝ث��_�61Nj48�.� H- �H�@R:_�L^ziPe��K�Я�F8\}�}�����Ћ� � Rk,�t�icMoj+@OoQxsp-@�"�3�CS jv+}LB-[5 HNj+� co~�L��z���f�k˝lb�jl!l����-˜�k/�.�x��LЎ�kipJ/�Gon,�J\A��8��SK"�� ��uto�o B������kwm� �o��H�tp�ʜ n}��exH-�˝��x���a^jIlL�je�식i���a��/���rej�1�o�V�or�zR����e qT�Z[��[lclN��߭�SOžGZD���to�{+B�H6343N�`�SG/o���sg�a�Utui��;`�J��`�;�;ndm�ndiN�{/ �/�/�/�/�/�/�/?`?/?A?�?��riΪ{! -Kj950/�sn �zk]895n/��O�t �Z��ws�g�K,�>��iag�� SGJ�Ю�o�gu���KO]Ltw�>_@	J64�1�sέ{F O>ګcdHݛ��`3_��r-�V�N74�y-�3��wRINnzlly���(m^���L���sg=c�zI" #?
+�oߡ\tw/��0�.�@�"���f�_�[yr�Kmm�K}dct^��t]�+�
PRZW7CHK
k,�;;`�y<p��lK���L.N*R85j �@_j�R ���tiN�g; WJhecN�L��F����wlZ|*��dat�ʛ�g�reN��o  �STD�r7LANG�Aoc�e�`��Q�y7��R870㕼{��8 (P�ogge���!��58\�PATT�s�� �t\��c "B�@V��1�Opatd���O����������{q㕔�5B�a�p[�m�\���7�\aw��@�a��p6�����ϯ�Ogmon���d� �0�B�m�;A��\ ö�K�I�MHCR��51 H����g�\o��@��R]� H#54ۿm�<@E���p;!�����omm�$;a��R�|�N㕬0�F�C��W�P�)Ai�6�� Fƫ�{��it�x�#{ ��iai�o����De6�ev9e����72 R�@tRƜPg��adl���nt��KRB�T�tOPTN�`772'�CTK�"'�g�(䔠�)� "AZ'�;q'�q'�'tzn&�{ E'�A{ma��- Mu���ncInDP�N�������87S2��|�d��(���������#���ma{sy��y "M��0o��䃲��et����\p1�����\ ��f���lZ����lp���9���`��+ V��ail��?��䇢�䄓���zd�<�k`��7�3.f��irdg.��- i��e\ ������ S0j�021"�1W ��(�`�4�n� (i��e,"�� "���+���coKre_�I��l`F��AY��AB��@�����H�����ABIC���Par;�M�ai�������<� c\ΖITX>���  {����1��wg Jclib��ShiW�4�� t�994\�VSS�F��� tt\j9�f "O�w� t��$%ini�/��pٰ t�5G�&,� t'\vsR&x�L�%w� tamclS/+rGef.�%#� tj�%m�� t[A�&4\9z�/�,z_v�%A8�%�a�%_ol6��8l% �%end�/<!c?.?@?R5o[?m>8�6�/�dshf�/+trt�?<OAE�'F  !�G��$%��Ƙ5vi�6���6 J�92�F3��%25 	(�%�@e&�P�%k�4O dnwzF��T�&`�XEpn�&g��?� nw\n�?�,n�d�V��N;XnF j���%se�V I/�
&�q&фU��5r w�%/F� �F�_�rclR&0\pw/Y��90�Eo`/"5�Of "U//A+dp�rm�%g¨%�Xrsu/kmS�T_ L`�6/OŔpM�LO�j��nO1|h�ODnon�|YCwrpR/�l���E�<�Pe\ga��Kr�gas�o�k��f�v��4xtf�?m$ra�o�la0�omk�_�TamN6+�4�`'9K0.v�Wې�%d�@�Ft��XE sV���ДJ737�%|�*�%,P��hB 9"+��KwcfF& �I����998�vt;omzFut vV�_�	o;�YC���:8\HF&�Y/� 0��f��deb^V��$�0�zFؠ"��g���<9)\�&��9�Wr}  �su"�st�G��X ؖf� U (�fag�n�F PzFϜ�Viaf�TX����vd���w��g��HzF- OƂW CH� �$723�F���E(A�ÿտ`2蚽Wc��WsvF&3 S�W�JR6��_�RVo RV���ӊ���vt�M\et(F�XoN�o�Fr��x����+�1T�F?teR�� J58�O  {34	Wgle,�%,�j�Dq\t"��zFfwIta1lUTA�VdϜ�gw韗Mad�Wp�Oa���6d M���e�FT��90 Hv�%NT��R69�ָ����ir\ʆM�IR��ӊenʆv���F|�3��ITCP���Ta0�p���(M�M7G�eT�o \t�pʆI��YBbusJ׈�m��I�@zFȀ���F�����/��W�'g, ��4`R_(!�sw�&s_YC67\JF��Tf_����D�fw��W��4ach�g��a96_��� _샏�_rV�%� 99YA�e���$FEAT�_ADD ?	������  	�$YA// %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�o�o# 5GYk}��� ������1�C� U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿�������DEMO N~�   �� *� �2�_�V�h��� ������������%�� .�[�R�d��������� ��������!*W N`������ ��&SJ\ �������� //"/O/F/X/�/|/ �/�/�/�/�/�/?? ?K?B?T?�?x?�?�? �?�?�?�?OOOGO >OPO}OtO�O�O�O�O �O�O___C_:_L_ y_p_�_�_�_�_�_�_ 	o oo?o6oHouolo ~o�o�o�o�o�o�o ;2Dqhz� ������
�7� .�@�m�d�v������� ƏЏ����3�*�<� i�`�r�������̟ ����/�&�8�e�\� n���������ȯ��� ��+�"�4�a�X�j��� ������Ŀ����'� �0�]�T�fϓϊϜ� ����������#��,� Y�P�bߏ߆ߘ߲߼� ��������(�U�L� ^���������� ����$�Q�H�Z��� ~�������������  MDV�z� �����
 I@Rv��� ���///E/</ N/{/r/�/�/�/�/�/ �/???A?8?J?w? n?�?�?�?�?�?�?O �?O=O4OFOsOjO|O �O�O�O�O�O_�O_ 9_0_B_o_f_x_�_�_ �_�_�_�_�_o5o,o >okoboto�o�o�o�o �o�o�o1(:g ^p������ � �-�$�6�c�Z�l� ��������Ə���� )� �2�_�V�h����� ��������%�� .�[�R�d�~������� ������!��*�W� N�`�z���������� ޿���&�S�J�\� vπϭϤ϶������� ��"�O�F�X�r�|� �ߠ߲��������� �K�B�T�n�x��� �����������G� >�P�j�t��������� ����C:L fp������ 	 ?6Hbl ������/� /;/2/D/^/h/�/�/ �/�/�/�/?�/
?7? .?@?Z?d?�?�?�?�? �?�?�?�?O3O*O<O VO`O�O�O�O�O�O�O �O�O_/_&_8_R_\_ �_�_�_�_�_�_�_�_ �_+o"o4oNoXo�o|o �o�o�o�o�o�o�o' 0JT�x�� �����#��,� F�P�}�t��������� ������(�B�L� y�p����������ܟ ���$�>�H�u�l� ~��������د�� � �:�D�q�h�z��� ����ݿԿ��
�� 6�@�m�d�vϣϚϬ� ���������2�<� i�`�rߟߖߨ����� �����.�8�e�\� n����������� ���*�4�a�X�j��� ������������ &0]Tf��� �����", YPb����� ���//(/U/L/ ^/�/�/�/�/�/�/�/ �/ ??$?Q?H?Z?�? ~?�?�?�?�?�?�?�? O OMODOVO�OzO�O �O�O�O�O�O�O__ I_@_R__v_�_�_�_�_�_�_m  h$o6oHoZolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ߀�߲����������  ��(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: L^p����� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p����� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺߠ��������� 	�,�>�P�b�t��� �����������(� :�L�^�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_��_�_�_�_oi�$�FEAT_DEM�OIN  d��D`�`,dINWDEX9kHa�,`�ILECOMP �O���za�Gb'ep`SET�UP2 Pze��b�  N ��amc_AP2BC�K 1Qzi G �)h�o�k%�o`}`Ae�o m�o� ��V� z�!��E��i�{� 
���.�ÏՏd����� ���*�S��w���� ��<�џ`������+� ��O�a�🅯���8� ��߯n����'�9�ȯ ]�쯁���"���F�ۿ �|�Ϡ�5�ĿB�k� ����ϳ���T���x� �߮�C���g�y�� ��,���P����߆�� ��?�Q���u���� :���^������)��� M���Z������6��� ��l���%7��[ ��� �D�h���i�`P�o }2�`*.VR`� *c�����JPC��� �FR6:�.�4/�TX`X/j/��U/�,;`%/�/�*#.FM�/�	��/�<�/<?�+STM@G?q?��]?�=+?�?�+H�?�?�7�?�?8�?EO�*GIFOOyO��5eO"O4O�O�*JPG�O�O�5�O�O�OM_F�JSW_�_� S�n_+_%
Java?Script�_�O�CS�_o�6�_�_ �%Cascad�ing Styl�e Sheets�0o� 
ARGNA�ME.DT_o��0\so1o�Q�d�o`o}�`DISP*�o �o�0�o7�e)q8�o�
TPEINS.gXMLg:\{�9�aCustom� Toolbar���iPASSWO�RD.�FRS�:\�� %P�assword ?Config@�� ���������r�� ���=�̏a�s���� &���J�\�񟀟��� �K�ڟo�������4� ɯX������#���G� ֯�}����0���׿ f������1���U�� yϋ�ϯ�>���b�t� 	ߘ�-߼�&�c��χ� ߽߫�L���p��� ��;���_��� ��$� ��H����~����7� I���m������2��� V���z���!��E�� >{
�.��d ��/�S�w �<�`�/ �+/�O/a/��// �/�/J/�/n/?�/�/ 9?�/]?�/V?�?"?�? F?�?�?|?O�?5OGO �?kO�?�OO0O�OTO �OxO�O_�OC_�Og_ y__�_,_�_�_b_�_ �_o�_�_Qo�_uoo no�o:o�o^o�o�o )�oM_�o�� 6H�l���7� �[����� ���D� ُ�z����3�ԏ i��������ßR�� v�����A�Пe�w� ���*���N�`���֦��$FILE_D�GBCK 1Q������� ( �)
�SUMMARY.�DG����MD:�3�s���Dia�g Summar�yt���
CONSLOGi�L�^��������Consol�e log����	?TPACCN�R��%:�wς�TP �Accounti�nρ�FR6:�IPKDMP.ZIP�ϯ�
���σ����Excepti�on ߱�_�MEMCHECKm�Կb�����Memor?y Data��֦�LN�)n�RI�PE�\�n����%�� Pack�et LϺ��$ySA���STAT������ߋ� %~�Status��<�	FTP����r������mmen�t TBD��� �=�)ETHERNEU���B�S������Ethern�(��figura�߇���DCSVRAF���������� verify �all٣M(=��DIFF�����/diff�PB���CHGD�1�x� X�FQ&��	28�� 5�YGD3���'/� �N/�UPDATES.m �S/��FRS:\�k/�-��Upda�tes List��/��PSRBWLOD.CM�/���"��/�/�PS_RO�BOWEL1���:GIG�ߊ?/�?�ֿGigE ��n�ostic*�ܢN��>�)�1HADOW�?�?�?5O���Shadow ?Change��٤�*8+�2NOT�I��O"O�O��N?otific��\O٥O�A��_�� 2_կ?_h_���__�_ �_Q_�_u_
oo�_@o �_dovoo�o)o�oMo �o�o�o�o<N�o r��7�[� ��&��J��W��� ���3�ȏڏi����� "�4�ÏX��|���� ��A�֟e�����0� ��T�f���������� O��s�����>�ͯ b��o���'���K�� 򿁿ϥ�:�L�ۿp� ���Ϧ�5���Y���}� ��$߳�H���l�~�� ��1�����g��ߋ� � 2���V���z�	��� ?���c���
���.���R�d�����������$FILE_� P�R� ����������M�DONLY 1Q����� 
 ��)�@_VDAEXTP.ZZZ���p�G�L6%N�O Back f�ile !��U3�M��7���� G�&�J\�� ��E�i�/ �4/�X/�e/�// �/A/�/�/w/?�/0? B?�/f?�/�?�?+?�? O?�?s?�?O�?>O�? bOtOO�O'O�O�O]O��O�O_(_��VIS�BCK����*�.VD)_s_�@F�R:\BPION\�DATA\^_R��@Vision VDt�_�O�_�_ _o_Ao�_Rowoo �o*o�o�o`o�o�o �o�oO�os�@� 8�\���'�� K�]�������4�F� ۏj����̏5�ďY� �j������B�ן� x����1���ҟg����MR2_GRP �1R���C4�  B�O�	 �
������E�� �֯�r���OHcE�P]��O��#�M��
�KA����?�&�r���:6:N�R��9-�Z��A��  v���BH��C`}dC��N��OB�{��r���xпὫ�@UUT���U����/Ϫ�>���>c��>r�а=ȫ�>�i�=���>�����:��:���:/:6?)�:��~ϗ� 2ϔ��ϸ������z�_CFG S��T  �a�s߅߾0[NO ���
F0�� ��/\R�M_CHKTYP  ���O�����������OM��_MsIN��L����v��X��SSB7�]T�� ���5�L�,�U�g���TP_DEF_OW���L�����IRCO�M�Ѝ��$GENOVRD_DO�ֹ	��THR�� �d��d��_ENB��� ��RAVCr��U�UQ �Υ m�X��|������n�� � �OU��-[��O�������8�:���x
,.  C��������h/�v%�������n�!�SMT'�\.���+��w�$HOSTC�7�1]K[��Y� 	MMdMI�}�e� ��� /*�1/C/�U/g/��/ 	anonymous�/ �/�/�/�/? L^ pM?�/� /�?�?�? �?/�?OO%O7OZ? �/�/O�O�O�O�O?  ?2?D?FO3_z?W_i_ {_�_�_�?�_�_�_�_ o._dOvOSoeowo�o �o�O�O_�ooN_ +=Oa�_r�� ���o�8o�'�9� K�]��o�o�o�o��� ����#�5�|Y� k�}�����ď��� ����1�x�����J� �������ӯ���	� ��-�?�Q�c�����Ο ����Ͽ��:�L�^� p�Mτ����ϕϧϹ� �������%�7�Z� ����ߑߣߵ����  �2�D�F�3�z�W�i� {������������� �
�d�A�S�e�w�����/ENT 1^��� P!���  ������* ��Nr5~Y� �����8� \1�U�y� ����4/�X// |/?/�/c/�/�/�/�/ �/?�/B??N?)?w? �?_?�?�?�?�?O�? ,O�?ObO%O�OIO�O�mJQUICC0 �O�O�O_�D1_�O�OV_�D2W_3_E_�_�!ROUTER�_�_�_�_!PC�JOG�_�_!�192.168.�0.10�O�CCA�MPRTGo#o!b7e1@`noUfRT�_�ro�o�o��NAME� !��!RO�BO`o�oS_CF�G 1]�� ��Auto�-started^��FTP��~q ���F����� ���9�K�]�o���� &���ɏۏ�����W i{X����o����� ğ֟������0�B� e��x���������ү �������Q�>���b� t�������q�ο�� ��9���L�^�pς� �Ϧ�������%�� Y�6�H�Z�l�3ϐߢ� ��������}��� �2� D�V�h���������� �����
��.�@�� d�v���������Q��� ��*<���� ��������� ���8J\n�� %�����EW i{}O/��/�/�/ �/�/��/??0?B? e/�/x?�?�?�?�?�? /+/=/�?Q?>O�/bO tO�O�O�Oq?�O�O�O _'O(_�OL_^_p_�_��_(�`_ERR �_z�_�VPDU�SIZ  9P^�S@��T>�UWR�D ?EuA� � guest3V$o6oHoZolo�~o�dSCD_GR�OUP 3`E| uIq?YM �nwCON�nTAS�n�L��nAXP�n_E��o9P�n�RTTP�_AUTH 1a��[ <!iPendan�g�~@}�9PJ�!KAR�EL:*���}�KC����pV�ISION SE!T�`E��I�!\�J� t��s����������Ώ���-���dtCTR/L b�]~�9Q�
@,FFF�9E39�DFR�S:DEFAUL�T��FANU�C Web Server����bvo dL��'�9�K�]�o��TWR_�`FIGw c�e�R����QIDL_C_PU_PC9QsB�@� BHǥ�MINҬ�a�GNR_IO�Q�R9P�X�ɠNPT_SIM�_DO�!�STAL_SCRN�� �y�+�TPMODNTOLY�!���RTY8��&�9�hp�ENBY��cƣO�LNK 1d�[ �`�����1�C�UϾͲMASTE����&�OSLAVE� e�_˴jqO_gCFGsϦ�UOD�|�Ϩ�CYCLE����ļ�_ASG 19f���Q
 W�9� K�]�o߁ߓߥ߷��߀�������#�_��N�UM�S�b�U
��I�PCH��j�O_R?TRY_CN�x�Z��U�_UPD�S����U �������g�θ`��`ɠP_�MEMBERS �2h��` $�e��>��HyɠSD�T_ISOLC � ���r�\J2/3_DS��q���?OBPROC��%��JOG�d1i���89Pd8�#?�.���.�?�?�?OQNs��V����3W~�����������POSR�E��$�KANJI�_m�K�i�pMO�N j�k~�9Ry ����//�^�r��k����9%Th���p_L�I�l�kEYLOGGIN����`����U�$�LANGUAGE� ����� ,�!�QLG��lq�9R마9Px�p�  ���砬9P'0�3X�k���MC�:\RSCH\0�0\��� N_DISP m��DA8MK�SLOCw�آ�Dz ��A�#OGBOOK nۄ��9P~��1�1�0X�9O%O7OIO[OmN`�Mɱ���I��	�5@Ib�5�O�O�5�2�_BUFF 1oؽ�O2A5!_�2 ��=_?7Y_k_�_�_�_ �_�_�_o�_o:o1o CoUogo�o�o�o�oe4~��DCS q�= =��͏L�O-��1CUg���bIOw 1r� ���s20����� ���1�A�S�e�y� ��������я���	���+�=�Q�|uE�TMl�d����Ο�� ���(�:�L�^�p� ��������ʯܯ� �8��7�SEV��u=]{�TYPl���`z�����!�PRS����/S��FL 1s�}����$�6�`H�Z�l�~ϯ�TP� �l�i��=NGNA�M��A5�"e4UPSFm0GI��\!�����_LOAD��G �%u:%REQ�MENU��3�MA?XUALRMI�c�8W�T���_PR�����3�R�Cp0t��9�M���3Eݗ���Pw 2u�� �1V�	i�00��� �߭�1��.�g�x U���������� ���8�J�-�n�Y��� u�����������" F1jM_�� �����	B %7xc���� ���/�/P/;/ t/_/�/�/�/�/�/�/ �/�/(??L?7?p?�? e?�?�?�?�?�? O�? $OOHOZO=O~OiO�O�K�D_LDXDI�SA����zsMEM�O_AP��E ?=��
 b��I �O_"_4_F_X_j_|_~R�ISC 1v�� ��O�_ ���_��_�Ooo@o�_C_MSTR w:�~_eSCD 1x�M�4o�o0o�o�o�o�o P;t_� �������� :�%�^�I���m���� ��܏Ǐ ��$��4� Z�E�~�i�����Ɵ�� �՟� ��D�/�h� S���w���¯���ѯ 
���.��R�=�O��� s�����п����߿� *��N�9�r�]ϖρ����PoMKCFG �ynm����LTAWRM_��z����и���6�>�s�M�ETPU�ӫІ��viND��ADCO�LXի�c�CMNT�y� l�g` {�nn��-�&�����l�P�OSCF����PgRPM����STw�{1|�[ 4@�P<#�
g��g�w� ��c��������� ����G�)�;�}�_��q�����������l�S�ING_CHK � |�$MODA�Q�}�σW��#D�EV 	�Z	�MC:WHSIZ�E�M�P�#TAS�K %�Z%$1�23456789� ��!TRIGW 1~�]l�U%�\�!�S
K.�S�Y�P�69"EM_INF 1�� `)�AT&FV0E�0X�)�E0�V1&A3&B1�&D2&S0&C�1S0=�)A#TZ�#/
$H'/O/�Cw/(A/�/b/�/�/�/? �&?� ��/�?3/�?�/�? �?�/�?�?"O4OOXO ??�OA?S?e?�O�? �?_CO0_�O�?f_!_ �_q_�_�_sO�_�O�O �O�O>o�Obo�_so�o K_�owo�o�o�o�_ �_L�_o#o��Yo ����o$��H� /�l�~�1��Ugy ���� �2�i�V�	��z�5�������ԟPN�ITOR��G ?�k   	EOXEC1���2�3�4�5�� �U7�8�9��� �������(���4��� @���L���X���d���Pp���|���2��2��U2��2��2��2ŨU2Ѩ2ݨ2�2���3��3��3(�#R�_GRP_SV �1�� (�ɳ�lC������6�MO�_Ds�����PL_NAME� !���!�Default� Persona�lity (from FD) ���RR2�� 1�L6(L?����	l d��nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ�������B2]��� *�<�N�`�r����<���������� ,�>�P�b�t�����B�J  ��\  �  ���Ȱ�  A� W B��T��� �
������� g ������B��p���  CH C�H P Ez � E�� E�` E�;%��Z�*� �  E��F[�@&��T Ai� dx�H �x�	$Hxd�
dڭ�}`( d��8(xx$$y Xtd D (DDdp WwX��	X�v@XHX���/yJ�y (� !���  7%E	��Em�Xw$%XH$%P�� �/�/�/�/ �/�/??+?=?O?a?s=F�r?�?�?�?��6��E�{PEWU���2 ��������?Kزd�� 'O9NO\OjG�0��|M���ز'4 � W%�O�O�N  �H�O�J�A  A��C�����_�OC_9W�  � TB�LY��
��_�\B��Q�Y=�CÈ��V�`HR0� ʒP( @7%?��a�Q�?ذaر@�6��&س��2n;�	l�b	  ����pX���U�M`�X� � � �,� �rb��K�l,�K���K��2�KI+�KG0�/K �U�L2o�E�	O�n��@6@� t�@�X@�I��b`�o�C��N����
���}v������` q�m�|�kQ�
=ô��  Hq�o~`!b���  Ȱ�a� ������ذa�s����}�m��o�q��v�O��E	'� � 0��I� �  �� Q�J:�È~T�È=���l���@|���}~�Q����R�����yN8���  '�<�ap?���b!p��b){�B��?�C�IpB  X��ذ���C�A�f��՚n`��(��BB P��8�����P��ԕرD �O���O���A�,���Š
��`l�1�	 S٠p��� p` l`�:GT  �t�?�ff{O��įV� �P�����a�!��/�?Y)R�a4�(ذ]�Pf����a\c\d^ƃ?333-d����;�x5;��0�;�i;�du;�t�<!�+}�oݯ��b�Sb�P�?fff?��?&���T@��A{#$�@�o[,� ��x�	�&f6�ed�g ���Hd㯸ϣ�����  ���$��H�Z�E�~���&eF��mߺ�i߀��U���y���2���E�0����y�d�� ������������ ?�*�܏r�8�.o�ߺ� ���T�);ڿ Pb��������P��A��T C�=�ϵ��Y}��2������m�C��W�C�= �` Ca��������(!�`�<����bC@_;C9��BA��Q�>V{È�����Y�?uü��
/�S���Q��hQ��A�B=�
�?h�Ä/iP�����W��ÈK��B/
=�����Ɗ=�K��=�J6XK��r#H�Y
H}���A�1�L��jLK����H:��H�K��/0	b�L �2J��8�H��H+UZBu�a?�/^? �?�?�?�?�?�?O�? O9O$O]OHO�OlO�O �O�O�O�O�O�O#__ G_2_k_V_{_�_�_�_ �_�_�_o�_1oo.o goRo�ovo�o�o�o�o �o	�o-Q<u `������� ��;�&�K�q�\���΀�Gϭ���� C�aɏ Ĉ�y���CVF������+b�����yKc�f�� 
E��Ў�T�ٟ��(���_3�h۟���������N�������3�lC�(�:�H�����T�f��t�.3礁}����k����q'�3�JJ �����گ���4�"�J]P̲Pf��������⟛�ſ���ԻA����/��?�{?�<N�u�  fUh�*� �Ϟ������Ϣ�t�.��R�@��X�bߘ�̆ߨ�)Z�ߺ�  ( 5�	�������B�0�f�t�  �2 E%p"E[[@��N�"B,C��%@ߏ��%��������;���������@����%n�n�%�đ�%��Xc
 ��!3EWi {��������b*[��P�I��v�$MSKCFMAP  ��� ^������pDONREoL  X�[���DEXCFEN�B�
Y�FN�C��JOGOV�LIM�d��d�DKEY��%_PAN�""�DRUN�+S?FSPDTYw��<��SIGN���T1MOT���D_CE_GRP� 1���[\ ���/��?&?��?Q? ?u?,?j?�?b?�?�? �?O�?)O;O�?_OO �O�OLO�OpO�O�O�O _%__I_ _m__f_��_O�DQZ_ED�IT�$UTCO�M_CFG 1�BQ�_o"o
�Q__ARC_�X���T_MN_MO�D���$�UA�P_CPLFo�N�OCHECK ?=Q W��� �o�o�o�o'9 K]o������vNO_WAITc_L�'�W� NT�Q��Q���_E�RR�!2�Q���� �_t��������*��Ώ�d``OI��>P�x Z�_�>��8�?0�4������B�PARAuMJ��Q���`	�����s�� =���345678901��� ���?�Q�-� ]�����u���ϯ����������7�ODRDSPEc�&��OFFSET_C�AR�PKom�DIS�z�K�PEN_FI�LE���!$a�V<`O�PTION_IO�
/!аM_PRGw %Q%$*	��ά�WORK ���'� ���K�7U�h��f�(�f�	 ���f�7����M�RG_D?SBL  Q������L�RIEN�TTO* ��C����Z��M�UT_S/IM_DطX+�M�VQ�LCT ��%��R_�$aQ�'�_�PEXh`��b�RA-Thg d�b�r��UP �5� �� ����߼������$��2�#�L6�(L?��	l d'�O�a�s�� ������������ '�9�K�]�o���������H�2>������/ASew�N�< �������@1CUgyH����P�� � � ��  �U�A��  B��PB�����H���  ���U�BJ�p������N��P Ez  E��� E�` EE��;(�����Z�/���  �E��''���@V#���T�AJ(��E!Y!a!)!m!Y!�u)%)!Y!E!�%E!��$�^$A!�	!E!a! �%%	-Y!Y%�-58��Z 99U%E!�D!	$D%%E!Q481X2 91�%�)95�/W#95)%�91m5a!�5/Z7��Z (�8�1�<a1 fEE	�(�Em�4�94X6E9=)%E15�� |O�O�O�O�O�O��O�O__0_B_T]F�S_y_�_�_�Vh������_�[��%� on�_=oKg�]�]&��'4 � �W%po�oX� �g��g�o�jA�A��c�����o�o$*w���tB�(~ �`��r�|�� q�y��$�O��1�+�k�+��3��`��0��P( @EhD�D��q?Q�C�Z7�}��o  ;�	l�D�	u� ���pX��[�2��X �� � �, ��W��`H��9H��H��H`��H^yH�R�l���_�����`�C#�B� C40ӄ����c�9��_�
=���� �������cBz���Βa�m�另b�s�� �q����g䟒�챏Ǒ��ٖ�o���e	'�� � �I� �  �q<�=���9�K���@a�g�b����������唠����N��  '۰��Ɓ"�B�Ղ��т6���� �  ���C�a����U��`��2�gBp ��Н����px����D��o޿�o��&�l�o�5�Ю`Q���	 ٠TU�f� U� Q�:����#����?�faf\o�ϩ�;� �p�����"�8� ��?%Y
r��q=�(� BՁPK�fɆ�A�A���?�333��m�;��x5;��0;��i;�du;�?t�<!��y�������t���r�p?f7ff?x�?&����@��A#	�@�o[�	]� �����uI��wh��� -��ϝ��������� 	���-�?�*�c�u�L� ������4�V�X����EjPf��^ I�m����  �$��W� ������9��/  /��5/G/�z/e/�/`�/�/�/�`�A��$�t�/ C�/"?�(���>�?��Pn?�/h�?}?��(��W�?{C�@�` CT���?�j4�j0i1A@�I�!���bC�@_;C9�B�A�Q�>�V`.È�����Y�uü��
�?�3��Q���hQ�A��B=�
?h���iOJp��W���ÈK�B/�
=�������=�=K�=�J�6XK�r#H��Y
H}��A��1�=L�j�LK����H:��HK���O�@	bL ��2J��8H���H+UZBu�?F_�OC_|_g_�_ �_�_�_�_�_�_o	o Bo-ofoQo�ouo�o�o �o�o�o�o,P ;`�q���� �����L�7�p� [��������ȏ�ُ ���6�!�Z�E�~�i� {�����؟ß��� ���0�V�A�z�e�G�y����� C�a�/>�� Ĉ��ЯׯOCVF�����üK<G�j���KH�K�� 
Ep�s�9���z90(91�_�h���y����i��N�����LA3lC�8��-¢�9�K���t�.3��}�e�w�k���q'�3�JJ�͑���@��������B5P��	PK�Zgt�ǿ��0�ߕ��߹�����߈���$�{$�3�Z�  fUM����� �����Y��7�%���=�G�}�k���)�Z����  ( 5�� ������'�KY  2 wE%pIFE[@t�N�IFB�!�!� C%��0� L@@į�����*H3 ��Tfx��LCLB94��L@D9=4H;
 �/ /*/</N/`/r/�/�/��/�/�/�/�/GJ@2���5�I�v�$�PARAM_ME�NU ?����  �DEFPULS���	WAITT�MOUTT;RC�Vg? SHE�LL_WRK.$�CUR_STYLv���<OPT�N�?PTB�?�2C�?R_DECSN_0 <�L	OO-OVOQOcO uO�O�O�O�O�O�O�O�_._)1SSREL?_ID  ��Y��=UUSE_PR_OG %8:%*_�_>SCCRk0ORY�@3�W_HOST !8:!�T�_�ZAT\Ю_ c�_�Qc|<o�[_TIMEi2�OV�U)0GDEB�UGMP8;>SGIN?P_FLMS`�gn�hTR�o�gPGA��` �lC�kCH��o�hTYPE5<A)_#_Y�}� �������� 1�Z�U�g�y������� ������	�2�-�?� Q�z�u�������ϟ��
��eWORD �?	8;
 	�PR�`��MAI�@��SU�1E�T1E#`���	�4R��COL��n���vT�RACECTL �1���B1 �I�W֯ࢵ�D/T Q����Р�D � ;��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� ����� $ 6@�bt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n�V���� ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z� �ߞ߰��ߘ����
� �.�@�R�d�v��� �����������*� <�N�`�r��������� ������&8J \n������ ��"4FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/?? ,?>?P?b?t?�?�?�?��?�?�?�?OC�$�PGTRACEL�EN  A  ��@��$F_UP �/���SA[@?A�  T@$A_CFG7 �SE=CAT@��D�D�O�G�6@�OhBDEFSP/D �sLA6@��$@H_CON?FIG �SE;CW @@dTM�3B AQP�DطA1Q@�$@IN~k@TRL �sM��A8�EFQPE�E�W�SA�DQ��ILIDlC�sM	~�TGRP 1�Y� lAC%�  ��l�AA��;H�N��R�A!PD	� a3C	\T�Ai�)iQP� 	 ��O4VGgCo ´|c^oGkB`�a�opo��o�o�o�o�b"�Bz�o7I~3� <}�<�oN�J���� �f�)��9�_�J�"`z����@
t��� d�ŏ�֏���3�� W�B�{�f�x�����՟������J)@)
�V7.10bet�a1�F @��@�A&�ff�Q2�CPC��`�D�Dk`[�C��T��@ DĠ� Dr� �QBH��`�L��PC5R �A?�  ��CCx����b��P!P��A,����Ap`B�bc0 ��$�6�eC�Q�KNOW_M  ��E{F�TSV �Z(R�C���� ��ʿ��ٿ�$�A�!m�SM�S�[ ��B�	�E��C�Ϗ�̓E`��2�E@�2������X��d@�QMR�S�Y�eT�j���ACf����e@�Rۚ]ST�Q1� 1�SK
 4 �U��,ժ߲C�ߡ߳� ��������-��1�v� U�g���������� ���	�N�-�?�Q�p��2{���A�<�����P3���������p�4��+p�5 HZl~p�6����p�7� $�p�8ASewp�M�AD0F [E��O�VLD  SK��ϼOr�PARNU�M  /]///T�_SCH� [E
�}'F!�)=C�%UPD�F/X%5U�/��_CM�P_O�0@T@@'�{E�$ER_CHK�5yH!6
?;RS8�]��Q_MO�o?�5_k?��_RES_GzФ~ݍ��?�O O�?%OO*O[ONOO rO�O�O�O�O�O�O��3���<�?_�5�� (_G_L_�3G g_�_�_ �3� �_�_�_�3� �_ o	o�3@$oCoHo�3��co�o�o�2V 1�~կ1e�@c?���2THR_IN�R�0�!7³5d�fM�ASS ZwM�N5sMON_QUEUE �~ըf��0���4N0U�H1NEv6;�pEND8�q�?�yEXE��u�� BE�p��sOP�TIO�w�;�pPR�OGRAM %�hz%�p�ol/�rT�ASK_I��~O?CFG �hZ/�\���DATARè.��@��2���� �#�5�G��k�}��� ����^�ן�������INFORé܍� wtȟe�w��������� ѯ�����+�=�O� a�s���������Ϳ(�4��܌ �I��� K_�����T��ENB� ͻ1>ƽ��I��G��2�� P(O�ҡϳ�� �����_E?DIT ����|ߋ�WERFL�x��cm�RGADJ {�8�A�  hՁ?�0t�
qLֈq����5�?��!��<@�x"*�%����@�#ߊ��2����F�	Hpl�G|�b��>��A�dw�t$I�*X�=/Z� **:c�0 V�h���Ǟ���B�����x"������� ������b���L�B� T���x���������: ����$,�Pb ������� ~(:h^p� �����V/ // @/6/H/�/l/~/�/�/ �/.?�/�/?? ?�? D?V?�?z?�?O�?�? �?�?�?rOO.O\ORO dO�O�O�O�O�O�OJ_ �O_4_*_<_�_`_r_ �_�_�_"o�_�_ooo�f	���o�p�o�o �dJ��oL��o#�oG�Y��PREF �����p�p
L�I�ORITY����>P�MPDSP�>�ƴwUTz�4�K�OD�UCTw�8��\�OG�_TG�;�|����rTOEN�T 1��� (�!AF_INE��pp�{�!tc�p{���!ud���ˎ!icmX�����rXY�Ӵ��;��q)� p�/�A��p�)�j�M�Y� ��}��������ן� ��8�J�1�n�U�����	*�s�Ӷ}}�����^,�>�%�jfp�!/z�֯K�,�������A��,  � �p�������ʿ�u"��ut�}�sF�P�PO�RT_NUM�s��p�P�_CARTREP�p��|��SKSTA�w nK�LGSm���������pUnothingϿ�������c{t�TEMP �����ke��_�a_seiban 0C�,S�y�dߝ߈� �߬�����	����?� *�c�N��r���� �������)��M�8� q�\�n����������� ����#I4mX �|�������3��VERSI��p �d disabled>SAVE ���	2600H7K21:&�!;�0��̏� 	(�r$moN+E/`�eb/�/�/�/�/�*z,�?� %`���_-� 1���E0�b8e�O?a?4gnpURGE_ENB3��v�u�WF�0DO�v��v�Wi��4�q*�WRU�P_DELAY ��CΡ5R_HOT %�f�q:�.O��5R_NORMA�LH
�OrOAGSE�MIQOwO�OlqQS�KIP-3���>3x $�O _1_C_]&o t_b_�_�_�_�_�_�_ �_o(o:o o^oLo�o �o�olo�o�o�o  $�oH6X~�� h��������D�2�h�z�����$�RBTIF�4G�R�CVTMOU\�v����DCR-3}��I �Q�/ Qʴ1Ed���A]	C����3=;4]�"�q&�j��QU��?�h�_�V�R_ ;�x5�;��0;�i�;�du;�t�<!��h��R���̝�����&�8� J�\�n�����������RDIO_TYP�E  4=��¯E�FPOS1 1�C�
 x/:�H2�� b�M���/��E�οi� ˿ϟ�(�ÿL��p� ���/�i��ϵ��ω� ߭�6���3�l�ߐ� +ߴ�O����߅ߗ��� 2��V���z���9� ����o�������@� R�����9���������OS2 1��; +�u���-��Q���3 1�����G����gS4 1�~���ZE~>�S5 1�%�7q��/�S6 1Ũ��/�/�o/�/&/S7 1� =/O/a/�/??=?�/S8 1��/�/�/�0?�?�?�?P?SMA_SK 1�߯ )�8OF�7XNOܯF�UO_C�MOTE��X4uA_CFG� �|M�1\A�P?L_RANGxA����AOWER ����@�FSM_D�RYPRG %��%y?!_�ETAR�T ��N/ZUME_PRO�O_�_�X4_EXEC_E�NB  ����GSPDdP�P�X���VgTDB�_�ZRM�_��XIA_OPTI�ONφ����pAI�NGVERS.a��z_�)I_�AIRPUR�@ q@O�o�=MT_�0�T�@zO��OBOT_ISOLC=N��F�1�a�eNA�MERl�bo�:OB�_ORD_NUM� ?�H�a�H721  �V1wLqr��qrV0qr��s�ps�u\@��PC_T�IMĖ��x��S7232�B1����a�LTEACH PENDAN΀��7\H��x?c��Maintena�nce Cons�V2�#�"�_�?No Use��N� �r���������С�rGNPO>P�r\A<e��qCH_LgP��|Nw�	<��!�UD1:b�	�R��0VAILRq2e���upASR  ��:a�B�R_�INTVAL1fᐄI�+n��V_D�ATA_GRP c2���qs0DҐP�?`��?��o���� ����կï����� -�/�A�w�e������� ���ѿ���=�+� a�Oυ�sϕϗϩ��� �����'��K�9�[� ��oߥߓ��߷����� �����G�5�k�Y�� }������������ 1��U�C�e�g�y��� ����������	+�Q?uDA�$SA�F_DO_PUL�S�pE@�C�� C�AN�r1f�vpS�C�@�+��+Ƙ�QV0D�D�qL�L�+AV2 y�'9 K]o��������ڈ���2($Md($C!8u�1#
) @�Co/ �/�/�.W)k/ M��$�_ @݃�T:`�/??&?39T D��3?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O֏<��i%�O�O��O܉�!L� �;��o݄�p�M
�?t��Dipp��L��J� � � �jL���j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������@���(�:����/ c�u���������Ϗ� �B�%�1�C�U�g� y���������Ƒ��0RMS�EW]�$�6� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ�����M�� �*�<�N�`�r߄ߖ� �����������&� 8�J�\�ǟ������� ������������,� >�P�b�p��������� ������%7I [m����� ��!3EWit�OB3t�� ���////A/S/ e/w/�/�/�/�/�/�*���/?6���\R?�M	12�345678XR�h!B!̺����?�? �?�?�?�?�?OOA �>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_o]-O�_�_�_�_ �_�_�_o"o4oFoXo�jo|o�o�o�oq_BH�o�o�o!3E Wi{���������v[;�j �A�S�e�w������� ��я�����+�=�O�a�xYD�k����� ��ɟ۟����#�5� G�Y�k�}�������v_ ׯ�����1�C�U� g�y���������ӿ� ��	�ȯ-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�σߕ� �߹���������%� 7�I�[�m�����"�v6����z���!�3�O:Cz  �A�z   ��@�2�v0� �@�
���  	�r������������Kph�u����� K]o����� ���#5GY k}��0��� �//1/C/U/g/y/ �/�/�/�/�/�/�/	?�?-?G�������*@ � <X4t��$SC�R_GRP 1��+� +�� �t �t�� E5	 /�1��2�2 �4��W1G3�;97�7�?8�?OC��|�B?D�` D��3�NGK)R-2�000iC/16�5F 56789�0��E��RC�65 �@�
1'234�E�6t�A�����C�1F�1 �3�1)�1A�:�1�I	��?_Q_c_u_�_~���H��0 T�7�2�_�?�_�_o�6�t��_Lo�_PpoB8boK�h�@��9�BǙ�B�  ?B�33Bƿ`�eȾb�c�1Ag��o  �@t��e�1@>@	 ' ?�w�bH�`2��j�1F@ F�`\rd[o�s�� �����*��k�c�)rU�@�R�d�v�B� ���ʏ���ُ��� �H�3�l�W���{����Ě2C�?���7����9�t�!q@"p6��G?�S�r�`y��`ȏ��G�L�3��ϯ�A>G�1��"o�e��)�t�  �<�N�\�*�q�}�\��^� P��(�����ӿ�g1EL_D�EFAULT  ��D���t���HOTST�R� ��MIPO�WERFL  �K����?�WFDO�� S�RVENT 1����P�0� L!DU�M_EIP翬���j!AF_IN�E��ϵ!FT$�������!�_B�� ��i�!RPC_MAINj��LغXߵ�|�VIS��Kٻ���!TMP��PU�߳�d���M�!
PMON_�PROXYN��e <���g��f�����!RDM_SR�V���g��1�!�R�DM���h �}�!%
~�M���il���!RLSYN�@�����8��!gROS��<�4�a!
CE�MT'COMb��kP�{!	vCONS����l��!vWOASRC ���m�vE!vUSBF��n4�0ߵ�� ��/�'/�K//�o/�RVICE_�KL ?%�� �(%SVCPR#G1v/�*�%2�/�/"� 3�/�/� 4??"� 56?;?� 6^?c?� 7�?�?� �D�?�,	9�?�;�$H�O�! �/+O�!�/SO�! ?{O �!(?�O�!P?�O�!x? �O�!�?_�!�?C_�! �?k_�!O�_�!AO�_ �!iO�_�!�Oo�!�O 3o�!�O[o�!	_�o�! 1_�o�!Y_�o�!�_�o �!�_{/�"� �/� F �E1������ ��
�C�U�@�y�d� ���������Џ��� �?�*�c�N���r��� �����̟��)�� M�8�_���n�����˯ ���گ�%��I�4� m�X���|�����ǿ��ֿρ*_DEV ����MC�:�H'�GRP� 2ׇ�+p� b�x 	� 
 ,y�ϒ�+r~ϻ� �����������9� � ]�o�Vߓ�z߷��߰� �����#�z�G���k� }�d���������� �����U�<�y�`� ��������*���	�� -QcJ�n� �����; "_FX����� ���/�/I/0/ m/T/�/�/�/�/�/�/ �/�/!??E?W?�{? 2?�?�?�?�?�?�?O �?/OOSO:OLO�OpO �O�O�O�O�O_^?�O =_�Oa_H_�_�_~_�_ �_�_�_�_o�_9oKo 2oooVo�ozo�o�o _ �o�o�o#
G.@ }d������ ��1��U�<�y��� �o��f�ӏ�̏	��� -�?�&�c�J���n��� �����ȟ����;� ��0�q�(���|���˯ ���֯�%��I�0� m��f�����ǿ����\��#�d ��	� 4��X�C�|�gϠϯ��%��������������������+� �O�=�s߁��Ϧ��� i����������	�� Q��x��A����� �������Y��P��� )���q����������� 1�U���I��Y m���	�-� !E3U{i� �����// A///Q/w/��/�g/ �/�/�/�/??=?/ d?v?-?O?)?�?�?�? �?�?OW?<O{?OoO ]OO�O�O�O�O�O/O _SO�OG_5_k_Y_{_ }_�_�__�_+_�_o oCo1ogoUowo�_�_ �oo�o�o�o	? -c�o��oS�O �����;�}b� �+���������ɏ� ݏ�U�:�y��m�[� �������ş�-�� Q�۟E�3�i�W���{� ���دꯡ�ï��� A�/�e�S���˯��� y��ѿ����=�+� aϣ���ǿQϻϩ��� �������9�{�`ߟ� )ߓ߁߷ߥ������� A�g�8�w��k�Y�� }��������=��� 1���A�g�U���y��� �������	��- =cQ������w ���)9_ ���O���� /�%/gL/^//7/ //�/�/�/�/�/?/ $?c/�/W?E?g?i?{? �?�?�??�?;?�?/O OSOAOcOeOwO�O�? �OO�O_�O+__O_ =___�O�O�_�O�_�_ �_o�_'ooKo�_ro �_;o�o7o�o�o�o�o �o#eoJ�o}k ������="� a�U�C�y�g����� ��ӏ���9�Ï-�� Q�?�u�c���ۏ��ҟ �������)��M�;� q�����ןa�˯��ۯ ݯ�%��I���p��� 9�����ǿ��׿ٿ� !�c�Hχ��{�iϟ� ���ϱ���)�O� �_� ��S�A�w�eߛ߉߿� ���%߯���)�O� =�s�a���߾��߇� ������%�K�9�o� �����_��������� ��!G��n��7 ������O 4F��g�� ���'/K�?/ -/O/Q/c/�/�/�/� �/#/�/??;?)?K? M?_?�?�/�?�/�?�? �?OO7O%OGO�?�? �O�?mO�O�O�O�O_ �O3_uOZ_�O#_�__ �_�_�_�_�_oM_2o q_�_eoSo�owo�o�o �o�o%o
Io�o=+ aO�s���o� !���9�'�]�K� �������q���m�ۏ ���5�#�Y������� I�����ßşן��� 1�s�X���!���y��� ������ӯ	�K�0�o� ��c�Q���u������� �7��G��;�)�_� Mσ�qϧ����ϗ� ߓ��7�%�[�I�� �Ϧ���o��������� �3�!�W��~��G� �����������	�/� q�V������w����� ������7�.�� ��O�s��� �3�'79K �o����� �#//3/5/G/}/� �/�m/�/�/�/�/? ?/?�/�/|?�/U?�? �?�?�?�?�?O]?BO �?OuOO�O�O�O�O �O�O5O_YO�OM_;_ q___�_�_�_�__�_ 1_�_%ooIo7omo[o }o�o�_�o	o�o�o�o !E3i�o�� Y{U����� A��h��1������� ��������[�@�� 	�s�a����������� �3��W��K�9�o� ]�����������/� ɯ#��G�5�k�Y��� ѯ������{���� �C�1�gϩ���ͿW� �ϯ��������	�?� ��fߥ�/ߙ߇߽߫� �������Y�>�}�� q�_�������� ��������7�m�[� ������������ ��!3iW��� ���}��� /e���U� ���/�/m� d/�=/�/�/�/�/�/ �/?E/*?i/�/]?�/ m?�?�?�?�?�??O A?�?5O#OYOGOiO�O }O�O�?�OO�O_�O 1__U_C_e_�_�O�_ �O{_�_�_	o�_-oo Qo�_xo�oAoco=o�o �o�o�o)koP�o �q����� �C(�g�[�I�� m�������ُ� �?� ɏ3�!�W�E�{�i��� ��؟������/� �S�A�w�����ݟg� ѯc�����+��O� ��v���?�����Ϳ�� ݿ��'�i�Nύ�� ��oϥϓ��Ϸ����� A�&�e���Y�G�}�k� �ߏ�������ߵ��� ���U�C�y�g����������$SER�V_MAIL  ������OU�TPUT����RV 2؍�  � (����_����SAVE���TOP10 2�9� d 	���� ����+=Oa s������� '9K]o� �������/ #/5/G/Y/k/}/�/�/��/���YP|���F�ZN_CFG �ڍ����j��!GRP 2���'&� ,B  � A=0��D;� �B>0�  B4~��RB21l�oHELL�"܍�$�L�M�7�?�;%RSR�?�?�?O �?%OOIO4OmOXOjO �O�O�O�O�O�O_!_~3^�  �R`3_a_s_AR_ ��1{_�R�P�xWIR�2��d�\�]�Rh6H�K 1�v;  �_o"ooFooojo|o �o�o�o�o�o�o�o�GBTfb<OM�M �v?�g2FTOV_ENB���A�$��ROW_RE�G_UI���IM�IOFWDL�p�x�~@5�WAIT�rA�Y�8���v@��0�TIM�u���j�VA��A��_U�NIT�s��$�LC��pTRY�w$����MON_ALI_AS ?e�yH�he��%�7�I�[�i� �������m���� 
��.�ٟR�d�v��� ��E���Я������ *�<�N�`��q����� ��̿w����&�8� �\�nπϒϤ�O��� ������߻�4�F�X� j�ߎߠ߲����߁� ����0�B���f�x� ����Y�������� ���>�P�b�t���� ����������( :L��p���� c�� �6H Zl~)���� ��/ /2/D/V// z/�/�/�/[/�/�/�/ 
??�/@?R?d?v?�? 3?�?�?�?�?�?�?O *O<ONO`OO�O�O�O �OeO�O�O__&_�O J_\_n_�_�_=_�_�_ �_�_�_�_"o4oFoXo oio�o�o�o�ooo�o �o0�oTfx ��G����� �,�>�P�b������ ����Ώy����(��:���$SMON�_DEFPRO ����c�� *S�YSTEM*M�R�ECALL ?}~c� ( �}A�@��şן���� �� 2�D�V�h�z������ ¯ԯ���
���.�@� R�d�v��������п ���ϙ�*�<�N�`� rτ�ϨϺ������� ߕ�&�8�J�\�n߀� ߤ߶��������ߑ߀"�4�F�X�j�|��}�+copy mc�:diocfgs�v.io md:�=>192.16�8.56.1:10496���������5��frs:o�rderfil.�dat virt:\temp\����g�y����-#�*.d7�I�Q�������xyzrate 61���������fx��8#�5�mpback��U��� }/��db��*���dv�6�3x�:\,��>YW��/�4�a��T�i/{/ �/��;V�/�/? �/B�/e?w?�?� //A/��?�?O/�? �?P/aOsO�O�/�/3? �/�O�O_?(?�OL? ]_o_�_�?�?9O�?�_ �_�_O$O�_HO�_ko}oo
# .o@oRo��o�o�#�D8220 �o�odv��o .@R���,16�p�� e�w����O�O7_8�ۏ ���_$_��7�ӏd� v����_,��o<�W�� ���o���p؟i� {�������;�V���� ����B�ԯe�w��� ��/�A�ҟ����� ����P�a�sυϘ��� 3�ί������(����L�]�o߁ߏ��$S�NPX_ASG �2�������  Z��%�����  ?����PARAM ����� �U	��P�������*����OFT_�KB_CFG  ��ô՞�OPIN_SIM  ��%�������RVQSTP_D�SBk�%����S�R �� �� &)�%�����T�OP_ON_ER�R  /�W�L�P_TN ����AH�RIN�G_PRMV� ���VCNT_GP� 2��'��x 	�������� ��$���VD��RP 1	���(���_ q������� %7I[m� �������/ !/3/Z/W/i/{/�/�/ �/�/�/�/�/ ??/? A?S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_r_o_ �_�_�_�_�_�_�_�_ o8o5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� ����	��-�?� Q�c�����������Ϗ ����)�P�M�_� q���������˟ݟ� ��%�7�I�[�m�� ������ܯٯ�����!�3�=PRG_CoOUNTL���[�_�ENB��Z�M���N䑿_UPD �1��T  
 H���ۿ���(�#�5� G�p�k�}Ϗϸϳ��� �� �����H�C�U� gߐߋߝ߯������� �� ��-�?�h�c�u� ������������ �@�;�M�_������� ����������% 7`[m��� ����83E W�{����� �/////X/S/e/ w/�/�/�/�/�/�/�/ ?0?+?=?O?x?s?�?�Q�_INFO 1Y�ɹ�� �F��?��?�?O�9���a�A��>>ܼO�;�S�Ɯ1���>O\�YSDEBSUGi�ʰ�0d���z@SP_PASS�i�B?�KLOG� �ɵ��r�0eH�?  �����1UD1:\x�DiO�A_MPC�M�ɵ:_L_ɱ�Aj_ �ɱVSAV �`�MA�A�B�5 X�SVnKTEM_T�IME 1��G.�� 0�0Y�4�U�oQ�T1SVGU�NSİj�'����`ASK_OPT�IONi�ɵ�����?a_DI�@��[eB�C2_GRP 2��ɹ�U�o�0@� � C��clBCC�FG �k�\ 9O
~`
EO B-Rxc��� ������>�)� b�M���q��������� ˏ��(��L�7�p����4m���n�ϟ� \�����;�&�_�q^ �QdT�������ѯ�� �����)�+�=�s� a���������߿Ϳ� ��9�'�]�Kρ�o� �ϓϥ����Ȭ���� �1�C���g�U�wߝ� �������߳�	���-� �Q�?�a�c�u��� ���������'�M� ;�q�_����������� ����7��Oa ��!���� �!3EiW� {�����/� ///S/A/w/e/�/�/ �/�/�/�/�/??)? +?=?s?a?�?M�?�? �?�?O�?'OO7O]O KO�O�O�OsO�O�O�O �O_�O!_#_5_k_Y_ �_}_�_�_�_�_�_o �_1ooUoCoyogo�o �o�o�o�o�o�?! ?Qc�o�u�� �����)��M� ;�q�_�������ˏ�� �ݏ��7�%�G�m� [��������ٟǟ� ���3�!�W�o��� ����ïA��կ��� �A�S�e�3���w��� ��ѿ������+�� O�=�s�aϗυϧ��� ��������9�'�I� K�]ߓ߁߷�m����� ���#��G�5�W�}� k����������� ��1��A�C�U���y� ������������- Q?uc��� ������/A _q�������/� �$TB�CSG_GRP �2����  �  
? ?�  J/\/ F/�/j/�/�/�/�/�/��/;#"*#�1,d�0?1?!	� HD 6@�Y3>��5O1B�H!x?�9D)��6L�ͣ1>���g6�0C�?�?�?�>p�?MCj���?5GB�B��OO)HY�0|Afff?IC�]O_O)O�2 �It?�N\0�/ XU&_ �O_Q_n_9_K_�_�_��[?��C �!�	�V3.00�R	�rc65�S	*`�T"o�V�4�T�p�Y G`mHo + � ��@�_�o��c#!J2*#�1-��o�hCFG ���;!C!�j�rB"]o~� BPz�Pva�� �������<� '�`�K���o������� ޏɏ��&��J�5� n�Y�k�����ȟ��� ���\	��-�ן`� K�p���������ޯɯ ��&�8��\�G��� k�����!/ۿ�� ���5�#�Y�G�}�k� �Ϗϱ���������� �C�1�S�U�gߝߋ� �߯�����	����?� -�c�Q���Y���� m������)��M�;� q�_������������� ����%I[m 9������� !E3iW�{ �����/�// /?/A/S/�/w/�/�/ �/�/�/�/?+?��C? U?g??�?�?�?�?�? �?�?OO9OKO]OoO -O�O�O�O�O�O�O�O _�O!_G_5_k_Y_�_ }_�_�_�_�_�_o�_ 1ooUoCoyogo�o�o �o�o�o�o�o	+ -?uc���� y?����;�)�_� M���q�������ݏ� ����7�%�[�I�� ������o�ٟǟ��� �3�!�W�E�{�i��� ������ï����� A�/�e�S�u������� ���ѿ�����+� a��yϋϝ�G��ϻ� �����'��K�9�o� �ߓߥ�c��߷����� ��#�5�G���}�k� ������������� �C�1�g�U���y��� ��������	��- Q?a�u��� ����/��� q_������ �/%/7/�/m/[/ �//�/�/�/�/�/? �/?!?3?i?W?�?{? �?�?�?�?�?O�?/O OSOAOwOeO�O�O�O �O�O�O�O__=_+_ M_s_a_�_C�_�_ }_�_�_o9o'o]oKo �ooo�o�o�o�o�o�o �o#Yk}� I������� ��U�C�y�g����� ����я����	�?� -�c�Q�s�u������� �ϟ��)�;��_S� e�w�!�����˯��ۯ ݯ�%��I�[�m���=�����ǿ���վ s �� ��)���$TBJO�P_GRP 2��ݵ� / ?��	A�H���O��� ����p{Xd� ���� � �,�� @�`�	 ߐD ��C?aD���`�x�¹���>���ϼ����<!a���?�����>L��?B�  B��8��C�D)�U�CQ?p�D�S�����>���u߻�ff�f���\<��Y�U��C +Р/�<��S�D5m�Κ��݁�&�)�333<���U�>���/>��C�й�<��b�Cj��u�b�����a�;�9b�B�!�?8Q��pG�Hc���s����Y��*��&�8��;��6��%�>u[%�DG���� ������*��8�&�<Z;u����� ����S�E/=k �w1����� ,�KeO]�d������ ��	V3.00f��rc65e�*� e��/ ' �F�  F�� �F� F�  �G� GX �G'� G;� �GR� Gj` �G�� G�| �G� G�� �G�8 G�� �G�< H� ?H� H��2 �Ez  E�@ _E�� EB F� �FR FZ F�� F� F�P<"G � GpL#�?h GV� G�nH G�� G��� G�( =^b�=+�8�$E�Q�?2�=3?�  ��M?�[:A��*SYS�TEM
!V8.3�0218 �38/�1/2017 �A y�p7M�T�P_THR_TA�BLE   $w $�1ENB��$DI_NO��O$DO�4���1�CFG_T � 0�0MAX_I�O_SCAN�2M;IN�2_TI�2D�ME\��0@�0 � � $C�OMMENT w$CVAL	C�T�0PT_IDXꉠEBL�0NUM�QBENDIJfAZIT�ID]B $D�UMMY13���$PS_OVERoFLOW�$�F��0FLA�0YP�E�2�BNC$GLB_TM�7�EF@�1��0ORQCTRL��1 X $DoEBUG�CRP�@�2@  $SB�R_PAM21_�VP T$SV�_ERR_MOD�U4SCL�@RAC�TIO�2�0GL_�VIEW�0 �4 $PA$Y*tRZtRWSPtR�A�$CA@A�1t�1aQUeU �0�N�P3@$GIF63@}$eQ lP_S��PiQ LpP�VI�<P�PF�RE�VNE�ARPLAN�A�$F	iDISTA�NCb�0JOG�_RADiQ�0$JOINTSPy尤TMSETiQ�  �WE�UAC�ONS2@B�RON�FiQ	� $�MOU1A`�$LOCK_FOL�A��2BGLV@CGL��hTEST_XM�@@raEMPE`,Rx�b�B`�$US;A�fPH`2P�S�aN�bMP_�`�aQ�CENEdRr $�KARE�@M�3T�PDRAhP;t2aV�ECLE�32dIU��aqHE�`TOcOLH`�0qsVI{s{RESpIS32�y;64�3ACHX`�`�~qONLE�D29��B�pI�1  �@$RAIL_B�OXEHaPRO�BO�d?�QHOWWAR�0�r�@�qOROLM�B�A�C� �SK�r�@�0O_F9�!��S�qiQ�
>o �RVpOC:iQ_�SLOGaK�[�UOUZbR��eAELECT�E<P`�$PIP�fNODE�r�r�q�IN�q2^��pCORDED�`�`}��0�P9P@  D� �@OBAU`T A�a����C�@���P8�q0��ADRA�0�F@TCHup � ,�0EN�2�1A
�a_�Tl�Z@�B�R�VWVA!A Ǥ ApeR�5PR�EV_RT�1$�EDIT��VSH�WR9�S@	UАIS|`yQ$IND0@�1QB蓗q$HEAD�5@ ��p5@���KEyQ�@CPSP]D�JMP�L�5��0RACE�4��a�It0S�CHANNEzp�	WOTICK{s�1M`Al�0@�HN�AD0Q^�]D�`CG�P����v�0STYf��qL�O�At����jP� t 
��Gr�%�$���T=PS�!$UNIGa5A�E��0�FPORT��SCQU5ptR���B��TERCJ@���T=SG� �PPL6�$�DE��$`Thqb�0OK@>CV�IZ�D4�Q�E�APR�A�Ͳ�1��PU}aݵ_�DObk�XSV`KN�6AXI��7�qgUR_s�E$T�p���*��0FREQ_,hp<�ET=�P�b�OPARA`@.P
@�:[���ATHr�3@a�D�s�s�0 ���SR_Q�0l8}��@�1TRQIc���$`�@��BRup��VyE@@��NOLD��AAp7a��x@�A��AV_MG����¨/���/�D)�D;�D�M�J_ACC.�C��<�CM��0CYC0M@3@��M@_E������٘@NbSSC��@  hPD1S���1�@SP�0*�AT:����@��i��B�ADDRES{sB���SHIF}b�a_%2��S@��I�@|�W�TV�bI�2]�гh>��C�
�j
#��V����0 \��������웱�@��CnӞ�aºꯆ:R����TXSCREE���0�TIN!AWS�P;��T�1>�>�jP TQ�7P�B �6QP��
��
�>��RROR_"a�@����D��UEG� ���U��@9SXQ�RSM�� �UNEXg��6��0S_�S��	0Ĭ�>�C�b��o� �26�UE����2GRUͰGMTN�_FLQ�#PO^HgBBL_�pWg@N�0 ����O�Q��LEn���pTyO`C�RIGH��BRDITd�CKG9Rg@�TEX,��>�WIDTH�sݐ�B�A�A{q �U�I_/@H�� 6� $LT_ �|�Y0@RyP�b�s�w�B��FOu��0D0$TW� U� �R�b��LUM�!�^�ERV��]PFP`>��1�'@r�GEUR��cF\��Q)��LP$�Z�Ed��)'��$(�$(�p#)5!+6
!+7!+8"b�>CȰP`��F�q�aS�@�EUSReT'  <��/@U�R��ξRFOChq�PPR�Iz�m�@?A� TR�IP�qm�UN�0�4!�P ��0�5��7��b;�5� "�T� ̱G �T07���}�O2OSNAd6ARA���;3wq�1#n_@�S�^�2����aU!"A$�?�?+"��;3�OFF�` P%O�z�3O@ 1#PtD,D$PGUN#�K`S�B_SUB8BPk SRT�0��a&��"avp��OR�pN�ERAU���DT�I�b��VCC��H�'� ��C36MF�B1ĢSPG?��( (b`�STEQʀ9PWTѠPEt���GXd) ����JMOVE��{Q6RAN4`?[�3DV�S6RLIM_X�3qV�3 qV\XvQk\:V1�IP�2VF��C���@d����*��IB�P,�S� _�`�p�b����@ (0G�B�� "P�@��pr+�x �r �,� tRn@��s C@TeGDRI�PSfQV!��wdԐ��D�$MY_UBY�$\d�;QA��S���h�q�bP_�S�ף�bL�BMvkQ$j�DEYg��EX� ���BUM_�MU6�X�D<q U�S��?��;VGo�PACI�TP�<Uyr��3yrkSyr:;qREnr�1l�8dyr�@�,�BTARGPP��q8eR{0�@- !d��;cB	:r���R�DSWqp�Sn�$:s˰O�!d�Av�3����E��U�p0m�V�vHK�.��K�`AQ��0���?SEA�����WOR�@3��uMwRCVr/ ��UO��M�@C�	Â8C�sÂREF�� ̆��gRj�
�� Ȋ��ي��=�̆r�_RC��s�����@������b�����A:bo0 ��Т�;��� �e�OU���r��\c(`	+�u��2��<���̰F� -=���f�K�WSUL3a.�C7Pfo/+p�NT�a ��]��ag��g��!g�&�L�c���c�����J�!�@T����1����o@AP_HU�R�ۥSA>SCMPB��F�����_&�AR�T������X.�ޗ�VGFS�E2d �M� � Y0UF_�����J���RO� ����W,rU�R�GR�mq�I ���D_V_h[D�@zYX��3�WIN.rH���X-V
A�RqR�P�WEw�w�q|c6v,q̓�RvLOiPtc��Ld��3t +�=�PA' =�CACH6����ŵ�,pP��2K�ۓC�QIo�FR"�T� $֭�$HO�@�R��`�rc ��[�֘p��ڔ��VP�r����_SZ�3p���6����12�� ��]p�؆P��WA�3�MP��aIMG�x���AD�qI�MREٔ6�_SI�Z�P��!po�6vA�SYNBUF6vV�RTDh�t�F�OLE_2D�T��t�J�0C0aUs��QP��X�ECCU�xVE�M�p����#�VIR9C��VTP������G�p��t��LA@�s�!��QMco4�0};�CKLASQCq	��ђ�@5  �AH�� @&B�T$��$`��6 |F@o���Xñ�T�o�?a��"¨uI���r/��`BGf� VEJ�`PK|pp1�1֖G�_HO+�>�R7 � }F�x��ESLOW}w�]RO>SACCE0*@-�=�xVR:��11�yrAD�/0r�PA��&�D�1��M_Ba�81��J�MP���A8y�b�O$SSC6u;�r)H��C��@92��S8�r��N/�PLEX��G: T〲C�Q��n6�FLD?1DEZ�FIQ rO�qty��F��PP2��;�� ϱPV多�MV_PIZ��G�BP0��`а�FIQ�PZ�$��������GA%p�LO9O0Tp�JCBT*����� ��ړPLAN�R&�L�F���cDV�'M�p���U�$�S�P.q�%�!�% #�㱶C4G�����RKE�1�VAN�C]G�A0p <��@�?�?J�R_A�a =�?q??T0�89��4�@> hܰ�	B��K9�fA2b<X@�̠OUe�ݒA��
�O���SK(�M�V{IE�p2= S08:�|R? <{@X�MԊ`UMMY��ԏ�Re��D��Ȧ�QCU�`b�U�@w@ $�@TIT 1�$PR8�UO�PT�VSHIyFʀ�A`�a`���T�0����$�_R$�UړQ.qZ� U�s�ot�Qav�Q�5fSTG@cVSCO��vQCNT���3�  }w�RlW�RzV�R�W�R��XLo^opjjA2���51D>a�0� .��SMO��B%X��J�@1u���_����@C%�Gi�L�I� '��XVR��DDY�@T�� Z7ABCP�E�r�btM��
�ZIP�EYF%��LV��L��z��bMPCF�eMGy�$p?�r?DMY_LN$@Aqq8��dH ����g��>�MCMİC>��CART_Xq��P�1 $JvsptD��|r�r�w��8�u���UXW�puUXEUL�x�q�u�t�u�q�q�y�q�vzZ�eI Hk��d���Y�`D�� �J 8o�	V�EgIGH��H?("��f��ĔK ��= �C���`$B&�Kģ��1_�B��LgRV� F^���COVC ؀qrfq9��@}�e��
����7�D�TR�Ȱ?�V�1�SPH� ǑL !�S�i�{�����ST�S  ����������u�<�ѐNa1 �� P������������U��������E��	���a������������������@��RDI�������ğ֟����t�O |���������ίஔ�	Sz��� >�����ſ ׿�����1�C�U� g�yϋϝϯ������� ���v�}���8�!�3� E�W���'�9�K�]�ؔ�� ��*��U��� A�@ ����0��@A�v�>^`BF_TT�������I�V>0n�J�_�I�R 1&�� 8����%к� ��C�  ������� �����"�4�F�X�j� |�������������1 gBTjx�����р��p��0B QI� ZlJ������ ���/"/4/F/X/ FҒ�t/�/b*���/�/���bv�@`�v�M�I_CHANU� "`� #3�dV�`�u��&0ET>�AD ?U��y0�m��/ �/�?�?�d0RLPs�!&�!�4�?�<?SNMASKn8���1255.4E0�33OEOWO�OOLOFS^Q �`�$X9�ORQCTRL &�V�m��O��T�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo(l�OKo:ooov��PE�pTAIL8��JPGL_CON?FIG 	�����/cell�/$CID$/grp1so�o�o1�#��?\n�� ��E����"� 4��X�j�|������� A�S������0�B� яf�x���������O� �����,�>�͟ߟ�t���������ίB�} c���(�:�L�^���`o��e��b���Ϳ߿ ���\�9�K�]�o� �ϓ�"Ϸ��������� �#߲�G�Y�k�}ߏ� ��0����������� ��C�U�g�y���� >�������	��-��� Q�c�u�������:��� ����);��_ q����H�� %7�[m�����]`��User Vie�w �i}}1234567890� 
//./@/R/Z$� �cz/���2�W�/ �/�/�/??u/�/�3�/d?v?�?�?�?�??�?�.4S?O*O<O@NO`OrO�?�O�.5O �O�O�O__&_�OG_�.6�O�_�_�_�_�_�_9_�_�.7o_4oFo�Xojo|o�o�_�o�.8 #o�o�o0B�o�cir l?Camera��o�������NE �,�>�P��j�|���0����ď�I  �v�) ��&�8�J�\�n�� �������ڟ����"�4�[��vR9˟�� ������ȯگ����� "�m�F�X�j�|����� G�Y�I7�����"� 4�F��j�|ώ�ٿ�� ��������߳�Y��� ��Z�l�~ߐߢߴ�[� ������G� �2�D�V� h�z�!߃unY����� ��������B�T�f� ��������������� Y�"i{�0BTfx �1����� ,>P��Y��i� �������/ ,/>/�b/t/�/�/�/�/cu9H/�/?!? 3?E?W?�h?�?�?F/ �?�?�?�?OO/O�j	�u0�?jO|O�O�O �O�Ok?�O�O_�?0_ B_T_f_x_�_1OCO�p �{._�_�_oo+o=o �Oaoso�o�_�o�o�o �o�o�_�u���oO as���Po�� �<�'�9�K�]�o� PEc����͏ߏ� ���9�K�]����� ������ɟ۟����ϻ r�'�9�K�]�o���(� ����ɯ�����#� 5�G��;�ޯ���� ��ɿۿ���#�5� ��Y�k�}Ϗϡϳ�Z� ����J����#�5�G� Y� �}ߏߡ����������������  ��N�`�r���������������   $�,�J�\�n��� �������������� "4FXj|�� �����0 BTfx���� ���//,/>/P/pb/t/�/�  
���(  �B�( 	 �/�/�/�/�/ ??8?&?H?J?\?�?��?�?�?�?�*4� �n�O1OCO��gO yO�O�O�O�O��O�O �O_VO3_E_W_i_{_ �_�O�_�_�__�_o o/oAoSo�_wo�o�o �_�o�o�o�o`o roOas�o��� ���8�'�9�� ]�o����������ۏ ���F�#�5�G�Y�k� }�ď֏��şן��� ��1�C�U���y��� �����ӯ���	�� b�?�Q�c��������� ��Ͽ�(�:��)�;� ��_�qσϕϧϹ� � �����H�%�7�I�[� m���ϣߵ������ ���!�3�E�ߞ�{� �������������� �d�A�S�e������ ��������*�+ r�Oas������0@ �������� ��)f�rh:\tpgl�\robots\r2000ic6�_165f.xml�`r����`���/����/ 3/E/W/i/{/�/�/�/ �/�/�/�//
?/?A? S?e?w?�?�?�?�?�? �?�??O+O=OOOaO sO�O�O�O�O�O�O�O O_'_9_K_]_o_�_ �_�_�_�_�_�__�_ #o5oGoYoko}o�o�o �o�o�o�o o�o1 CUgy���� ���o��-�?�Q� c�u���������Ϗ�t�K �� 88�?� �2��.�P�R�d��� �������П��� (�R�<�^���r������ܫ�$TPGL_�OUTPUT ����� ����%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{Ϡ�ϟϱ�����ˠ2�345678901��������0�8� ����_�q߃ߕߧ߹� Q߽�����%�7���}A�i�{����I� [�������/�A��� O�w���������W��� ��+=����s �����e� '9K�Y�� ���as�/#/ 5/G/Y/�g/�/�/�/ �/�/o/�/??1?C? U?�/�/�?�?�?�?�? �?}?�?O-O?OQOcO �?qO�O�O�O�O�OyO֡}�_)_;_M___�q_�]@��_�_�? ( 	 ���_ �_o�_5o#oYoGoio ko}o�o�o�o�o�o�o /UCyg� �������	�?��Ƭ�-�G�u��� c�������ߏ���`� �,�ΏP�b�@����� ���Οp�ޟ���� :�L���p���$����� ��ܯ�X���$�Ư� Z�l�J������ƿؿ z�����2�DϮ�0� zό�.ϰ��Ϡ����� b��.���R�d�B�t� �������߄��� ��<�N��r��&�� �������Z�l�&�8� ��\�n�L�������� ��|����� FX ��|�0���� �d0� fx V�����/ /�>/P/�</�/�/�:/�/�/�/�/?
2��$TPOFF_L�IM [��@W����A2N_S]V#0  �T5:�P_MON �S�74�@�@2��U1STRTCHOK S�56_�=2VTCOMPA�TJ8�196VWVA/R j=�8N4� �? O�@�}21_DEFP�ROG %�:%�&OmO;4_DISP�LAY*0�>?BIN�ST_MSK  �L {JINU�SER�?�DLCK��L�KQUICKM�EN�O�DSCRE�PS��2tpsc�D�A1P6Y52�GP_KYST�:59R�ACE_CFG ��Fr1�4.0	�D
?��XHNL 2�93��Q�; $B�_�_o o2oDo�Vohozj�UITEM� 2�[ �%�$1234567�890�o�e  =�<�o�o�os  !{!@�oZC �o{�o���9 K�o/��?�e�� ����#���G�� �+���O���ŏ׏Q� ����͟ߟC��g�y� ���]����������� �-���Q��u�5�G� ��]�ϯ!����ſ)� տ���q�ϕ����� 3�ݿ�ϯ���%���I� [�m���	ߣ�c�u��� �������3���W�� )��?���ߌ��ߧ� ����c�S�e�w�� �����k�������� +�=�O���s�EW ��c������9 �o��n� ����#�G� "/}=/�M/s/�/� �///1/�/U/?'? 9?�/]?�/�/�/i?�? ?�?�?Q?�?u?�?PO �?kO�?�O�OO�O)O(;O_�TS�R�_UJ��  �bUJq �Q`_UI
 m_�_z_�_8ZUD1�:\�\��QR_�GRP 1�k� 	 @`@ o!koAo/oeoSo�own��`�o�j�a�_�ox�o�e?�  ' 9{#YG}k�� �������C�`1�g�U�w���	�E���ÏSSCB 2%[ �!� 3�E�W�i�{�����\�V_CONFIG %]�Q]_�_����OUTPUT �%Y���� �S�e�w��������� ѯ�����+�_A@� S�e�w���������ѿ �����+�<�O�a� sυϗϩϻ������� ��'�8�K�]�o߁� �ߥ߷���������� #�5�F�Y�k�}��� ������������1� B�U�g�y��������� ������	->�Q cu������ �);L_q �������/ /%/7/H[/m//�/ �/�/�/�/�/�/?!? 3?D/W?i?{?�?�?�? �?�?�?�?OO/OAO ݟ�>�O�O�O�O�O �O�O�O_!_3_E_W_ J?{_�_�_�_�_�_�_ �_oo/oAoSod_wo �o�o�o�o�o�o�o +=Oaro�� �������'� 9�K�]�n�������� ɏۏ����#�5�G� Y�j�}�������şן �����1�C�U�g� x���������ӯ��� 	��-�?�Q�c�t��� ������Ͽ���� )�;�M�_�p��ϕϧ� ����������%�7� I�[�m�~ϑߣߵ��� �������!�3�E�W�|i�LH����� ���s���hO����� �1�C�U�g�y����� ����t�����	- ?Qcu���� ����);M _q������ �//%/7/I/[/m/ /�/�/�/�/��/�/ ?!?3?E?W?i?{?�? �?�?�?�?�/�?OO /OAOSOeOwO�O�O�O �O�O�?�O__+_=_ O_a_s_�_�_�_�_�_ �O�_oo'o9oKo]o oo�o�o�o�o�o�o�_ �o#5GYk} ������o�� �1�C�U�g�y��������ӏ���$TX�_SCREEN �1�����}��&�8�J�\�n��������� ҟ���������P� b�t�������!�ίE� ���(�:�L�ïp� 篔�����ʿܿ�e� w�$�6�H�Z�l�~��� ������������ � ��D߻�h�zߌߞ߰� ��9�K���
��.�@� R���v��ߚ����������k���$UA�LRM_MSG k?��� � �zJ�\����������� ��������/"SF|w+�SEV  ��E��)�ECFoG ���  �u@�  }A�   B��t
 x�s� 0BTfx�������GRP 2�� 0�v	 ��/+�I_BB�L_NOTE ��
T��#l�r��q� +"�DEFPRO5�%9� (%k�/�p �/�/�/�/�/?�/%? ?6?[?F??j?�?!,�INUSER  �o-/�?I_MENHIST 18���  (� � ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1�?`OrO�OΖO�� (O:M936MO�O�O__�B/_ A_S_e_w_�_�_*_�_ �_�_�_oo�_=oOo aoso�o�o&o�o�o�o �o'�oK]o ���4���� �#��<V""A�_�q� ���������ݏ�� �%�7�Ə[�m���� ����D�V�����!� 3�E�ԟi�{������� ïR������/�A� Я�w���������ѿ `�����+�=�O�:� L��ϗϩϻ������ ��'�9�K�]��ρ� �ߥ߷�������|�� #�5�G�Y�k��ߏ�� ��������x���1� C�U�g�y�������� ��������-?Q cu`�rϫ��� �);M_q ������/ /�7/I/[/m//�/  /�/�/�/�/�/?�/ 3?E?W?i?{?�?�?.? �?�?�?�?OO�?AO SOeOwO�O�O���O �O�O__+_.OO_a_ s_�_�_�_8_J_�_�_ oo'o9o�_]ooo�o �o�o�oFo�o�o�o #5�o�ok}�� ��T����1� C��g�y�����������O��$UI_P�ANEDATA �1������  	�}ӏ�,�>�P�b�t� )v���V��şן �������C�*�g� y�`������������ ޯ��?�Q�8�u�R�� �A������ Ŀֿ����_�0ϣ� B�f�xϊϜϮ���'� ��������>�%�b� I߆ߘ�߼ߣ�������7���T�Y� k�}�������J� ����1�C�U���y� ��r�����������	 ��-QcJ�n ��0�B��) ;M�q���� ���/h%//I/ 0/m//f/�/�/�/�/ �/�/�/!?3??W?� ��?�?�?�?�?�?:? OO�AOSOeOwO�O �OO�O�O�O�O�O_  _=_O_6_s_Z_�_�_ �_�_�_�_d?v?4O9o Ko]ooo�o�o�_�o*O �o�o�o#5�oY kR�v���� ���1�C�*�g�N� ����o"oӏ���	� �-���Q��ou����� ����ϟ�H���)� �M�_�F���j����� ��ݯį����7��� ��m��������ǿ� ���p�!�3�E�W�i� {�⿟φ����ϼ��� ���/��S�:�w߉��p߭ߔ���D�V�}�����-�?�Q�c�u�) 	��ŉ��������� � ���D�+�h�O�a� �������������� @R9v	�`�Z���$UI_POSTYPE  `��� 	 ����QUICKMEN  ����� REST�ORE 1 `��  �	i�S`N�m~������ /%/7/I/[/�/�/ �/�/�/r�/�/�/j/ 3?E?W?i?{??�?�? �?�?�?�?�?O/OAO SOeO?rO�O�OO�O �O�O__�O=_O_a_ s_�_(_�_�_�_�_�_ �O�_o"o�_Fooo�o �o�o�oZo�o�o�o #�oGYk}�:o ���2���1� C��g�y����������d����	��-��S�CRE� ?��u1scH�u2h�3h�4h�5*h�6h�7h�8h���USERJ�O�a�TLI�j�ksr�є4єU5є6є7є8ё�� NDO_CFG� !����Ѩ P�DATE ����None �_� ��_INFO� 1"`�]�0%3�x�	�f�����˯ ݯ������7��[� m�P�������ǿ�J��OFFSET %�ԿσA֏� *�<�N�{�rτϱϨ� ��Ͼ����A�8� J�w�n߀ߒ������
����UFRA_ME  ʄ��G�RTOL_AB�RT&��>�ENB�G�8�GRP 1&�<Cz  A�����������@������:�� Ug���V�MSK  (j�]�X�N#���]��%�߫��VCCMf�'���RG��E*�	��ʄƉ]D � BH)�p<�2C�)��PN?ـ` ��MR��20���p���"�р	 ����~XC56 �*������N�5р�A@<C�� ��� ʈ);h�c�"�Rр|��Ђ B��� �6�t/T1/ / U/@/y/d/�/�/�/�/ */�/	?�/???�c?\u?��TCC��1��Pf�9�рр��GFS�22w� Й�2345678901�?�2ʈ "�6��?!Oс>,12�$QO_GB@R 8N?:�o=L�� ���������OO A�O�O@O_dOvO�O �O�O�_�O�O�___ �_<_N_`_r_Soeo�_ Ro�o�_�_oo&o8o|��4SELECF��j�$�VIR�TSYNC� ���6�BqSIONT�MOU-tр���cu��3U���U�(�� �FR:\es\+�A�\�o �� �MC�vLOG� �  UD1�vE�X�с' B�@ ����q�DESKTOP-?8U37T7F�6���q:�^�σ ��  =	 1-� n6  -��ʆ�xf,p�#�0O=��ʹ���r}�xTRAIN�P�2�1.��
. d��t�sq4w (,1 ��0��)�;�M�_�q� ��������˟ݟ����I��crSTAT' 5��@�o��ĩ�E:$��ۯ�_GuE��6w�`. ��
��. 2�HO�MIN��7U��U� �r�a�a��aCG�um�JMPERR 28w
  ʯE:��su Ts�����߿��� '�9�O�]ώρϓ�_v-_�pRE��9t����LEX��:wA1�-e�VMPHA�SE  RuCCb��OFFLpc�<v�P2�t;4�04��8���b@�� �b<b>?s33��Á�1��L��ҕԈ�|��t�>x��Â�xf��o.���/?P�X� $�2�x����0�  ���6�+���l�� \�j�|����������  �D�V���ZTf ����������.  �,BPb�� �����// (/:/�y/�b/��/ �/L/? ??<?n/ c?�/�/�?�?�/�?6? �?�?�?OX?j?\O�? �OJO�?fO�O�O�O�O 0O%_TO_xOm_�O�O �O�_�_�_�__o>_ P_EoWo�_xo�_�o�o��o�o��TD_FI�LTEt�?�� ��Wp��]o$6 HZl~���� ����)�;�M��_�q������SHI�FTMENU 1-@x�<��%��� ��я��0���f�=� O���s�����䟻�͟����P�'�	L�IVE/SNAP�D�vsfliv��b���IO�N G�U���menu����:������l����A���	�����b�K��5M����m`@�����A�pB8������Ӝѝ�r�����m`� ;�,��/�ME��uYѵ�M���MO��B����z��WAIT�DINEND��3���OKN�.�O�UT#��Sa�4�T�IM�����G Ϯ�@���`ϱ�ϱ����2�RELEAS1E����TM���{��_ACTx���Ȫ�2�_DATA' C�ի�%i���<����RDIS�b޿�$XVR2�D���$ZABC_�GRP 1E8��n`,@h2��ǽZIP1�FD� cCo�������x�MPCF_G' 1G8�n`0<o ����=�H8����t�� 	�w�  8�R�����e�����?�k������5��
�\��  �a ������7�����I��z��Y�LIND�aJ��� �f ,(  *s�K�p���� �//+. mN/�r/Y/k/�/� �/�/�/3/?�/�/J? 1?n?U?�/�?�?v�C�s2K8��� �� O`o�7O~[Ol�?��Og��AA�AS�PHERE 2LS�?�OX?�O__ >_�?�Ot_�_?�_I_ /_�_�_o�_]_:oLo �_�_�o�_�o�o�o�o`#o $7�ZZ� �k�