��   �A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ��
��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !  �FTP_CTRL.� @� LOG_�8	�CMO>$�DNLD_FIL�TER�SUBD_IRCAP� �HO��NT. �4� H�9ADDORTYP� A H� �NGTHOG���z +LS/ D� $ROBOTyIG BPEER�ބ MASK@MR�U~OMGDEV�K���RCM+?� :$�� ���QSIZNT�IM$STA�TUS_�?MA�ILSERV�  �$PLANT� <�$LIN�<$C�LU��f<$TO�cP$CC5&FR\5&JEC!��ENB � ALkAR�B�TP��w#�V8 S��$�VAR)M�ONxt&��t&APPLt&�PA� u%�s'PO�R �_T!["AL�ERT5&2URL� }�#ATT�AC[0ERR_oTHRO�#US29�38� CH- �[4wMAX?WS_1w�y1MOD�z1I� $y2 � }(y1PWD  ; cLAu00�NDq1�TRY�6DELA��3z0��1ERSI�S�!�2�RO�9C�LK�8M� ��0X�ML+ �#SGFR�M�#TCP�OU��#PING_RE�5OP�!UF�#[A�qC�"u%_B_AUZ�@��B�!DUMM�Y1��A2?P_�RDM*�_$DIS�"� {SM� l5��!,"%�'NICC"b%H � 0VR#01U�P*_DLVP+AR��J@Io/ }3 $ARP��)_IPFOW_x��F_IN�FAD� �HO�_� INFO��wTELs	 P~���� WOR~�1$ACCE� �LV�[�"�I�CE�0 a  ��$�S  ��)�@a��
��
5`P�SlA>g%5�PbI0AL=oOaX'0 ^h
���F��a��%�b�e��� �m��!Ga�o����$ETH_FL�TR  ]i�` U��������{��� �m2{�RSH�cPD 1�i G P�o��d� ������:�� F�!�o���W���{�܏ �� �Ï$����Z�� ~�A���e�Ɵ������ �� ��D��h�+�a� ����¯��毩�
�ͯ ��?�d�'���K��� o�п������ɿ*�� N��r�5ϖ�Y�k��� ���ϳ����8���1߀n�]ߒ�U߶�wz _�L�11}x!�1.��0��y���1|�y�255.9�L����ܶe��2�߀�m��.�@�R�d�3 n����������d�4���]���0�B�d�5^��������������6���M ��� 2����6A�MY� MY����p{�K`�� Q� ��~< �/SewJ��v�P���/ �%/7/I/[///�/�/~t/uٹe�/�,��/i/2?D?V?h?}�}�iRConnect: irc�4�//alerts m?�?�?�?�?x5,?O@#O5OGOYOkO}��c9d�`pd��pO�O �O�O�O�O __$_6_ H_Z_l_~_{�$ O�_`p(�_�_$?�_oo�+oy�:`p�� �\b�jNeKabe|�Suֿ DM�c�n�$�SMIu�{��%�_�o�$`p�o}���o8#\�,��TCWPIP�b�m�(,�~qEL��	�eSa��  H!T�Phs�rj3�_tp�Bp|��Pq!KCL��{P|��>f!CRT@��.�����!C�ONS���z�qs'mon���