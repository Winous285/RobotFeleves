��   ��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A 	  ����DRYRUN_�T   � }$'ENB 4 �NUM_PORT�A ESU@$STATE P _TCOL_��PM�PMCmGRP_�MASKZE� O�TIONNLOG�_INFONiA�VcFLTR_E�MPTYd $P�ROD__ L �E�STOP_DSB�LAPOW_REwCOVAOPR��SAW_� G %$INIT	�RESUME_T�YPEN &J_�  4 $�($FST_ID1X�P_ICI0 �MIX_BG-yA
_NAMc �MODc_US�d�IFY_TI� xMKR�-  $L{INc   �_SIZcv� k�. , $USE_FL4 �p�&i*SIMA��Q#QB6'SC�AN�AXS+IN�S*I��_COUN�rRO��_!_TMR_VA�g�h>�i) �'�` ��R��!�+W[AR�$}H�!�{#NPCH���$$CLASS ? ���01���5��5%0VERS��.7  ��
A1IRTU�� .?@0'/ l5W5��������Y0�6m071�5��%@71�?���?
O��}5I2�;�GOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_���%FW?N8�0 ���_J�[m0�]��o { 2�;G 4%t_$o���1 �1oWo6o{o�olo�o�o�o�o��8�o���G" 
O��= q">���" wry@�S���=�9Y0��1�t�1�tX�1l1 Y0�>�&�8�J�\�n� ��������ȏڏ��� �6�1��1 �2�D�V� h�z�������ԟ����
�44�6�S!2>�9 �[� m��������ǯٯ� ���!�3� �M�f�x� ��������ҿ���� �,�>�I�b�tφϘ� �ϼ���������(� :�L�W�p߂ߔߦ߸� ������ ��$�6�H� S�e�~�������� ����� �2�D�V�a� z��������������� 
.@Rdo�� ������ *<N`k}�� ����//&/8/ J/\/n/�V