��   m�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����DMR_GRP�_T  � �$MA��R_D�ONE  $�OT_MINUS�   	GPyLN8COUNP �T REF>wP�OOtlTpB�CKLSH_SI�GoSEACHMsST>pSPC�
��MOVB RAD�APT_INERzP �FRIC�
_COL_P M�
�GRAV��� HsIS��DSP?��HIFT_ER[RO�  �NA�pMCHY SwARM_PARA#w d7ANGC �M2pCLDE|�CALIB� �DB$GEARz�2� RING���<$1_8k�  �FMS*�t *v M_LIF��u,(8*���M(DSTB0+_0>*_���*#z&~+CL_TIM��PCCOMi�F�Bk M� �MAL�_�EC�S�P�!Q%XO g$PS� �TI����%�"r $DT�Y?R. l*1EN�D14�$1�ACT�1#4V22\93\94�\95\96\6_OVR\6� GA[7�2h7 �2u7�2�7�2�7�2�8oFRMZ\6DE�{DX\6CURL� 
HSZ27Fh1DGu1�DG�1DG�1DG�1DCN�A!1?( �P�L� + ��S�TA23TRQ_Mȫ�/@K"�FSX��JY�JZ�II�JI��JI�D �$U1S�S  ����6Q����+PVE�RSI� 4W� �
GQIRT�UAL3_EQ' 1� TX  
��(P���_�_�_ �_o�_%oo"o[oFj� zjco?S�o�o �$7@�v����������-� �o�o�o�l/VSe�k��r�������d�#�5�<G���=L��R�y�3?�z���@����� я�����+�=�O�0a�s���� rU��p����ޟ:T  2� �!�3�E�W�i�{���������<��ۯ��� �#�5�G�Y�k�}��������sP��$$ �1�\�qKb��L��K���E�� N׿��N(���}J���wKb)0K�Dy6!�E8��D#���}o@�}�1�}�� ZϘ�Wϐ�{ϴ�'�9� �����.��R�=�v߈� ��ߓ�t���������UBu+UPz�q�6���Z� l�~�=�O������� ��� �2���V�h�z� 9�K�����������
 .��Rdv5G �����* �N`r1C�� ���//&/�J/ \/n/-/?/�/�/�/�/ �/�/?"?���/J?\? n?�/�?�?�?�?�?�? �?O"O�?FOXOjO)O �O�O�O�O�O�O�O_�_�OB_T_f_��,(�$1234567890�_�U���_�_ �_�_�_�_oo;o+o GoOoao�o�o�o�o�o �o�o�oI9U ]y������ �!��-�5�G�{�k��������ՏŅ�$P�LCLų�� Dm�?�  �1�%�T� m�x�c����������� �����>�P�