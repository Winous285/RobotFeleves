��   b�A��*SYST�EM*��V8.3�0218 8/�1/2017 �A   ����CELLSET�_T   �w$GI_STY�SEL_P }7T  7ISO:iRibDiTRA�R�>�I_INI; �����bU9AR�TaRSRPNS�1Q234�5678�Q
TROBQACKSNO� �)�7�E�S �a�o�zU2 3 4 5 6 7 8awn&GINm'D�&��) %��)4%��)P%�̖)l%SN�{(OU���!7� OPTNAA�73�73.:B<;�}a6.:C<;CK;C�aI_DECSN�A�3R�3�TRY�1��4��4�PTHCN�8D�D�INCYC@HG��KD�TASKOK �{D�{D�7:�E� U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V�8�Tb@SEGq�Tp��T�@REQ� d�drG�:Mf�GJO_HFAUL�Xpd�dvgALE�  �g�c�g�cvgE� �H<�dvgNDBR�H�dgRGAB�Xtb�  �CLML�Iy@   �$TYPESI�NDEXS�$$�CLASS  ���lq��;pup�apVERSION�ix  ��
}qIRTUAALi{q'61�r���p��q�t+ U�P0 �xS�tyle Select 	  ����r�uReq. /�Echo���A�ck���Initiat�p�r�E
�^�m����ʠ�	��
��  ���������������χ�q)��O�ption biGt A<��p�B���C4�Decis��codY��Tr?yout mj�6��Path seg�h�ntin.8�I�g�ycX�:�Tas�k OK��?�Ma�nual optK.r�A���B����C� decs�n ��$�Robo�t interl�o7�@�\� iso)lQ�4�C��iM�@���ment<�)��������Ě}�stat�us=�	MH F�ault:����Aler�1�C��p@r7 1�z j�;��y���I�; LE_COMNT ?�y�   Չ�ѿ �����*�<�N�`� rυϖϨϺ������� ��&�9�J�\�n߀� �ߤ߶����������"�����U��Ђ��Ŵ�   ��ENAB  ��:��������������ꮵME�NU\��y��NAM�E ?%��(%$*R�זb��P���t� ��������������+ O:s^p�� ���� $ 6HZ�~��� ����/ /Y/D/ }/h/�/�/�/�/�/�/ �/?
?C?.?@?R?d? v?�?�?�?�?�?�?�? OM