��   ��A��*SYST�EM*��V8.3�0218 8/�1/2017 �A 	  ����PASSNAM�E_T   0� $+ �$'WORD  �? LEVEL � $TI- OU�TT  &F/�� $SET�UPJPROGR�AMJINSTA�LLJY  ?$CURR_O��USER�NUM��STPS_LOkG_P N��$�eT�N�  6 �COUNT_DO�WN�$ENB�_PCMPWD �� DV�IN�!$C� CR=E�PARM:� =T:DIAG:)|�LVCHK!>FULLM0��YXT�CNTD��MENU�A�UTO,�FG_wDSP�RLS��U�fENC/�  CRY�PTE   �  �$$CL�(   ����;!�� D 0 V� I�O� :& � �
L!IRT�UA� :/�$DC�S_COD@�|��?%�  W�'�_S  v*�!$x �&�A91�"w!�� 
 $ B!���-�/? ?6?D? Z?h?~?�?�?�?�?�?��?�?OO2O���#SUP� �+4OFO�#�FfOxO�O��B, �L�A���O � ��� V�[t�&��j���D �ON_��W
_��d �V�x_UCLUGH 1}w) d �)�_�_�_oo)o ;oMo_oqo�o�o�o�' �_�o�o�o/A Sew����o� ����+�=�O�a� s���������ߏ� ��'�9�K�]�o��� ������Ə۟���� #�5�G�Y�k�}����� ��¯�����1� C�U�g�y��������� Я���	��-�?�Q� c�uχϙϫϽ�̿�� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ������������!� 3�E�W�i�{������� ��������/A Sew����� �%